DTLG �         @0����Name|Group|Class  @0����Units @0����Description 
@SData  � �       CalVIEW - RT Types.ctl g@ U8U32I8I32SGL	TBL1D_SGL	TBL2D_SGLU32_ENUMBOOLArray1D_SGLArray2D_SGLSTRCalVIEW Types @!Control  P          @ ����                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   :   'DrivvenReserved|Reserved|Target_Version       CalVIEW Target Version �                       )DrivvenReserved|Reserved|Protocol_Version       CalVIEW Protocol Version �                       #DrivvenReserved|Reserved|IP_Address       Target IP Address �     0����      
10.15.1.55            DrivvenReserved|Reserved|OS_Name       Target OS Name �     0����      PharLap           #DrivvenReserved|Reserved|OS_Version       Target OS Version �     0����      13.1            DrivvenReserved|Reserved|App_Env   finvalid app kind|Development System|Run Time System|Student Edition|Embedded LabVIEW|Evaluation|Custom   Target Application Environment �                       #DrivvenReserved|Reserved|Target_CPU   \invalid CPU target|Motorola 68K|PowerPC|Intel x86|SPARC|PA-RISC|MIPS|Alpha|ARM|AMD/Intel x64   Target CPU Type �                       "DrivvenReserved|Reserved|Target_OS   �invalid OS target|Mac OS|Windows 3.1|Windows 95/NT|Solaris 1|Solaris 2|HP-UX|PowerMAX|Linux|Irix|Rhapsody|BeOS|AIX|OSF1|VxWorks|PharLap|Carbon|RTX|Windows x64|Linux x64   Target OS Type �                       )DrivvenReserved|Reserved|Default_Data_Dir       Target Default Data Directory �     0����      c:\ni-rt\LabVIEW Data            DrivvenReserved|Reserved|IO_Lock   LOCKED|UNLOCKED   I/O Hardware Lock �     !               "DrivvenReserved|Reserved|Host_Time       Host Computer Timestamp �         �!�#           $DrivvenReserved|Reserved|Target_Time       Target Timestamp �         �!a�           *DrivvenReserved|Reserved|CalFile_Save_Time       Last Calibration File Save Time �     0����      13:16:55 08/02/2013           $DrivvenReserved|Reserved|Target_Name       Target Machine Name �     0����      NI-PXI8108-2F14CA16           "DrivvenReserved|Reserved|Host_Name       Host Machine Name �     0����      NILT-S7R160OZC0           %DrivvenReserved|Reserved|CalFile_Name       Calibration File Name �     0����      
DefaultCal           $DrivvenReserved|Reserved|Free_Memory   MB   -For Internal Use Only - Free Memory on Target �     	    ��             "DrivvenReserved|Reserved|Free_Disk   MB   Free Disk Space on Target �     	    ��              DrivvenReserved|Reserved|CPU_Use   %    For Internal Use Only - CPU Load �     	    ��             &DrivvenReserved|Reserved|CalVIEW_Build       CalVIEW Build Number �     0����      3.120.10700           $DrivvenReserved|Reserved|Scope_Count       For Internal Use Only �                      %DrivvenReserved|Reserved|Scope_Memory       For Internal Use Only �     	   @ ����                                              	    (DrivvenReserved|Reserved|Scope_Control_0       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_1       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_2       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_3       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_4       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_5       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_6       For Internal Use Only �     	   @ ����               	    (DrivvenReserved|Reserved|Scope_Control_7       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_0       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_1       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_2       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_3       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_4       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_5       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_6       For Internal Use Only �     	   @ ����               	    %DrivvenReserved|Reserved|Scope_Data_7       For Internal Use Only �     	   @ ����               	    .DrivvenReserved|Reserved|Non_Atomic_Array_Read       For Internal Use Only �                        /DrivvenReserved|Reserved|Non_Atomic_String_Read       For Internal Use Only �                        "DrivvenReserved|Reserved|IO_Locked   LOCKED|UNLOCKED   For Internal Use Only �     !               DCAT|AO|AO Type       2Analog output type associate with the measurement. �     	   @ ����               	   DCAT|AO|Cylinder       *Cylinder associated with each measurement. �     	   @ ����               	   DCAT|AO|Disable       LDisables data acquisition and calculations associated with each measurement. �     	   @ ����               	   DCAT|AO|Gain       &Gain associated with each measurement. �     	   @ ����               	   DCAT|AO|Max       5Maximum voltage range associate with the measurement. �     	   @ ����               	   DCAT|AO|Min       5Minimum voltage range associate with the measurement. �     	   @ ����               	   DCAT|AO|Name       5Name or description associated with each measurement. �     0����                 DCAT|AO|Offset       (Offset associated with each measurement. �     	   @ ����               	   DCAT|AO|Physical Channel       2Physical channel associated with each measurement. �     0����                 DCAT|AO|Type       2Measurement Type associated with each measurement. �     	   @ ����               	   DCAT|Async Digital|Cylinder       9Cylinders associated with each measurement in a bitfield. �     	   @ ����       G� G� G� G�                                                        	   DCAT|Async Digital|Invert       <Invert the digital signals associated with each measurement. �     	   @ ����                                                                              	   DCAT|Async Digital|Name       &Name associated with each measurement. �     0����      gTDC;Data;Reduce Resolution;Reserved;DI 4;DI 5;DI 6;DI 7;DI 8;DI 9;DI 10;DI 11;DI 12;DI 13;DI 14;DI 15
          DCAT|Async Digital|Type       2Measurement Type associated with each measurement. �     	   @ ����                                                                              	   DCAT|Async|Cylinder       9Cylinders associated with each measurement in a bitfield. �     	   @ ����               	   DCAT|Async|Disable       LDisables data acquisition and calculations associated with each measurement. �     	   @ ����               	   DCAT|Async|Filter       HFilter resource number associated with each measurement. (0 = No Filter) �     	   @ ����               	   DCAT|Async|Gain       cGain associated with each measurement when using  the gain only or gain and offset scaling methods. �     	   @ ����               	   DCAT|Async|Max       ?Maximum channel voltage range associated with each measurement. �     	   @ ����               	   DCAT|Async|Min       ?Minimum channel voltage range associated with each measurement. �     	   @ ����               	   DCAT|Async|Name       5Name or description associated with each measurement. �     0����                 DCAT|Async|Offset       VOffset associated with each measurement when using the gain and offset scaling method. �     	   @ ����               	   DCAT|Async|Physical Channel       2Physical channel associated with each measurement. �     0����                 "DCAT|Async|Polynomial Coefficients       bPolynomial Coefficients associated with each measurement when using the polynomial scaling method. �     	   @ ��������                         
   DCAT|Async|Scaling       0Scaling method associated with each measurement. �     	   @ ����               	   DCAT|Async|Table X       STable X array associated with each measurement when using the table scaling method. �     	   @ ��������                         
   DCAT|Async|Table Y       STable Y array associated with each measurement when using the table scaling method. �     	   @ ��������                         
   !DCAT|Async|Terminal Configuration       >Terminal Configuration array associated with each measurement. �     	   @ ����               	   DCAT|Async|Type       2Measurement Type associated with each measurement. �     	   @ ����               	   DCAT|Async|Units       'Units associated with each measurement. �     0����                 DCAT|Basic|Endpoint Window   CAD   iSpecifies the size of the window used to average the endpoints when calculating the polytropic exponents. �     	    @             DCAT|Basic|Exhaust Pressure End   CAD   6Specifies the end of the exhaust pressure calculation. �     	    C�            !DCAT|Basic|Exhaust Pressure Start   CAD   8Specifies the start of the exhaust pressure calculation. �     	    C�            DCAT|Basic|Intake Pressure End   CAD   5Specifies the end of the intake pressure calculation. �     	    Ö             DCAT|Basic|Intake Pressure Start   CAD   7Specifies the start of the intake pressure calculation. �     	    ô            DCAT|Basic|Peak Pressure   Standard|Spline (Very Slow)   9Specifies the method used to calculate the peak pressure. �                       DCAT|Basic|Peak Pressure End   CAD   .Specifies the end of the peak pressure window. �     	    Bp            DCAT|Basic|Peak Pressure Start   CAD   0Specifies the start of the peak pressure window. �     	    �p            DCAT|Basic|Polytropic   !Point-byPoint|Endpoints|Power Fit   @Specifies the method used to calculate the polytropic exponents. �                       %DCAT|Basic|Polytropic Compression End   CAD   <Specifies the end of the polytropic compression calculation. �     	    �p            'DCAT|Basic|Polytropic Compression Start   CAD   >Specifies the start of the polytropic compression calculation. �     	    ´            #DCAT|Basic|Polytropic Expansion End   CAD   :Specifies the end of the polytropic expansion calculation. �     	    B�            %DCAT|Basic|Polytropic Expansion Start   CAD   <Specifies the start of the polytropic expansion calculation. �     	    Bp            DCAT|Buffer|Alignment Overflow   	Overflow|   'Indicates an Alignment buffer overflow. �     !               DCAT|Buffer|Alignment Queue   %   #Indicates the Alignment buffer use. �     	                   DCAT|Buffer|Async Ind Overflow   	Overflow|   ;Indicates an overflow of Asynchronous Index process buffer. �     !               !DCAT|Buffer|Async Ind Process Use   %   4Indicates the Asynchronous Index process buffer use. �     	                   "DCAT|Buffer|Async Ind Raw Overflow   |   <Indicates an overflow of Asynchronous Index raw file buffer. �     !               %DCAT|Buffer|Async Ind Raw Process Use   %   5Indicates the Asynchronous Index raw file buffer use. �     	                   DCAT|Buffer|Async Ind Raw Use       5Indicates the Asynchronous Index raw file buffer use. �                        DCAT|Buffer|Async Ind Size       4Indicates the size of the Asynchronous Index buffer. �                        DCAT|Buffer|Async Ind Use       4Indicates the Asynchronous Index process buffer use. �                        DCAT|Buffer|Async Overflow   	Overflow|   5Indicates an overflow of Asynchronous process buffer. �     !               DCAT|Buffer|Async Process Use   %   .Indicates the Asynchronous process buffer use. �     	                   DCAT|Buffer|Async Raw Overflow   |   6Indicates an overflow of Asynchronous raw file buffer. �     !               !DCAT|Buffer|Async Raw Process Use   %   /Indicates the Asynchronous raw file buffer use. �     	                   DCAT|Buffer|Async Raw Use       /Indicates the Asynchronous raw file buffer use. �                        DCAT|Buffer|Async Size       .Indicates the size of the Asynchronous buffer. �                        DCAT|Buffer|Async Use       .Indicates the Asynchronous process buffer use. �                        DCAT|Buffer|Cycle Data Overflow   	Overflow|   'Indicates a Cycle Data buffer overflow. �     !               DCAT|Buffer|Cycle Data Queue   %   $Indicates the Cycle Data buffer use. �     	                   DCAT|Buffer|Display Overflow   	Overflow|   $Indicates a Display buffer overflow. �     !               DCAT|Buffer|Display Queue   %   !Indicates the Display buffer use. �     	                   DCAT|Buffer|FPGA Overflow   	Overflow|   -Indicates an overflow of FPGA process buffer. �     !               DCAT|Buffer|FPGA Process Use   %   &Indicates the FPGA process buffer use. �     	                   DCAT|Buffer|FPGA Raw Overflow   |   .Indicates an overflow of FPGA raw file buffer. �     !                DCAT|Buffer|FPGA Raw Process Use   %   'Indicates the FPGA raw file buffer use. �     	                   DCAT|Buffer|FPGA Raw Use       'Indicates the FPGA raw file buffer use. �                        DCAT|Buffer|FPGA Size       &Indicates the size of the FPGA buffer. �                        DCAT|Buffer|FPGA Use       &Indicates the FPGA process buffer use. �                        DCAT|Buffer|Feedback Overflow   	Overflow|   %Indicates a Feedback buffer overflow. �     !               DCAT|Buffer|Feedback Queue   %   "Indicates the Feedback buffer use. �     	                   !DCAT|Buffer|Medium Speed Overflow   	Overflow|   5Indicates an overflow of Medium Speed process buffer. �     !               $DCAT|Buffer|Medium Speed Process Use   %   .Indicates the Medium Speed process buffer use. �     	                   %DCAT|Buffer|Medium Speed Raw Overflow   |   6Indicates an overflow of Medium Speed raw file buffer. �     !               (DCAT|Buffer|Medium Speed Raw Process Use   %   /Indicates the Medium Speed raw file buffer use. �     	                    DCAT|Buffer|Medium Speed Raw Use       /Indicates the Medium Speed raw file buffer use. �                        DCAT|Buffer|Medium Speed Size       .Indicates the size of the Medium Speed buffer. �                        DCAT|Buffer|Medium Speed Use       .Indicates the Medium Speed process buffer use. �                        DCAT|Buffer|Next-Cycle Ready   CAD   ]Indicates the crank angle where the Next Cycle Data became ready for use in the control loop. �     	                   DCAT|Buffer|Raw File Overflow   	Overflow|   %Indicates a Raw File buffer overflow. �     !               DCAT|Buffer|Raw File Queue   %   "Indicates the Raw File buffer use. �     	                   !DCAT|Buffer|Summary File Overflow   	Overflow|   )Indicates a Summary File buffer overflow. �     !               DCAT|Buffer|Summary File Queue   %   &Indicates the Summary File buffer use. �     	                   DCAT|Buffer|Sync Overflow   	Overflow|   4Indicates an overflow of Synchronous process buffer. �     !               DCAT|Buffer|Sync Process Use   %   -Indicates the Synchronous process buffer use. �     	                   DCAT|Buffer|Sync Raw Overflow   |   5Indicates an overflow of Synchronous raw file buffer. �     !                DCAT|Buffer|Sync Raw Process Use   %   .Indicates the Synchronous raw file buffer use. �     	                   DCAT|Buffer|Sync Raw Use       .Indicates the Synchronous raw file buffer use. �                        DCAT|Buffer|Sync Size       -Indicates the size of the Synchronous buffer. �                        DCAT|Buffer|Sync Use       -Indicates the Synchronous process buffer use. �                        DCAT|Calculations|Basic   Enabled|Disabled   Enables the Basic calculations. �     !             DCAT|Calculations|Cam   Enabled|Disabled   Enables the Cam calculations. �     !              DCAT|Calculations|FPGA   Enabled|Disabled   Enables the FPGA calculations. �     !              DCAT|Calculations|Gas Temp   Enabled|Disabled   )Enables the Gas Temperature calculations. �     !              DCAT|Calculations|Heat Release   Enabled|Disabled   &Enables the Heat Release calculations. �     !              DCAT|Calculations|Injector   Enabled|Disabled   "Enables the Injector calculations. �     !              DCAT|Calculations|Knock   Enabled|Disabled   Enables the Knock calculations. �     !              DCAT|Calculations|MEP   Enabled|Disabled   1Enables the Mean Effective Pressure calculations. �     !              DCAT|Calculations|Medium Speed   Enabled|Disabled   1Enables the Mean Effective Pressure calculations. �     !             DCAT|Calculations|Misfire   Enabled|Disabled   !Enables the Misfire calculations. �     !              DCAT|Calculations|Motoring   Enabled|Disabled   "Enables the Motoring calculations. �     !              DCAT|Calculations|Noise   Enabled|Disabled   Enables the Noise calculations. �     !              DCAT|Calculations|PWM   Enabled|Disabled   0Enables the Pulse Width Modulation calculations. �     !              DCAT|Calculations|Pump   Enabled|Disabled   *Enables the Synchronous Pump calculations. �     !              DCAT|Calculations|Spark   Enabled|Disabled   Enables the Spark calculations. �     !              #DCAT|Calculations|User Calculations   Enabled|Disabled   Enables the User calculations. �     !              #DCAT|Calculations|User Heat Release   Enabled|Disabled   3Indicates whether the user heat release is enabled. �     !               DCAT|Calculations|User Process   Enabled|Disabled   Enables the User Processing. �     !               DCAT|Cam|Exhaust Cam Edge Angles   CAD   @Specifies the angle for each exhaust cam pulse of each cylinder. �     	   @ ��������                                                                                                                                                                                                                                                                                                                                                                                                                 
   DCAT|Cam|Exhaust Cam Edge Count       =Specifies the number of exhaust cam pulses for each cylinder. �     	   @ ����                                                                              	   $DCAT|Cam|Exhaust Cam Edge Directions   CAD   �Specifies the direction of exhaust cam pulse for each cylinder. Each cylinders data is stored in a bit field corresponding to each pulse. �     	   @ ����                                                                              	   DCAT|Cam|Intake Cam Edge Angles   CAD   >Specifies the angle for each input cam pulse of each cylinder. �     	   @ ��������                                                                                                                                                                                                                                                                                                                                                                                                                 
   DCAT|Cam|Intake Cam Edge Count       <Specifies the number of intake cam pulses for each cylinder. �     	   @ ����                                                                              	   #DCAT|Cam|Intake Cam Edge Directions       �Specifies the direction of intake cam pulse for each cylinder. Each cylinders data is stored in a bit field corresponding to each pulse. �     	   @ ����                                                                              	   DCAT|Control|Buffer Size   s   *Specifies the minimum size of the buffers. �     	    ?�            DCAT|Control|Current Units       "Specifies a list of current units. �     0����      kPa;kPa abs;ns;kW          DCAT|Control|Desired Units       "Specifies a list of desired units. �     0����      psi;psia;sec;hp          DCAT|Control|EPT Sim Enable   Simulation|Engine   EEnables EPT simulation of engine encoder signals for offline testing. �     !              DCAT|Control|EPT Sim Speed   RPM   +Setpoint for simulated EPT encoder signals. �     	    Dz            $DCAT|Control|Enable Unit Conversions   Enabled|Disabled   *Enables unit conversions on host displays. �     !              DCAT|Control|Knock Period   ms   &Specifies the update rate on host VIs. �           �          DCAT|Control|Next-Cycle Cutoff   CAD   USpecifies the angle to process Next-Cycle data. Any data after the cutoff is invalid. �     	    Bp            DCAT|Control|Next-Cycle Enable   Enabled|Disabled   ?Enables Next-Cycle calculations for the engine controller code. �     !             DCAT|Control|Plot End   CAD   JMaximum crank angle to display on a plot when using a custom global scale. �     	    C�            DCAT|Control|Plot Period   ms   &Specifies the update rate on host VIs. �            d          DCAT|Control|Plot Scale   \No Change|Autoscale|Custom|-360 to +360|-180 to +180|-60 to +60|-30 to +30|0 to +60|0 to +30   <Global control of all plots with Crank Angle for the X-Axis. �                      DCAT|Control|Plot Start   to   JMinimum crank angle to display on a plot when using a custom global scale. �     	    ô            DCAT|Control|Pre-Triggered Size   Cycles   -Specifies the number of pre-triggered cycles. �            
          DCAT|Control|Rolling Stats Size       5Specifies the size of the rolling statistics buffers. �            d          DCAT|Control|Run State   	Setup|Run   8Controls the state of the DCAT DAQ tasks and processing. �     !             #DCAT|Control|Save Trigger Direction   Rising|Falling   2Specifies the direction for the save file trigger. �                       #DCAT|Control|Save Trigger Threshold       5Specifies the threshold used for a save file trigger. �     	    ?�            DCAT|Control|Simulation   Enabled|Disabled   3Enables a simulation that doesn't require hardware. �     !              DCAT|Control|Start Delay   ms   &Specifies the start delay of host VIs. �           �          $DCAT|Control|Statistics Refresh Rate   ms   &Specifies the statistics refresh rate. �            d          DCAT|Control|Table Period   ms   &Specifies the update rate on host VIs. �            d          DCAT|Control|Trend Period   ms   &Specifies the update rate on host VIs. �           �          DCAT|Control|Trigger Size   Cycles   1Specifies the number of cycles to save at a time. �            
          DCAT|Control|Unit Multiplier       SSpecifies the conversion factor to get from the current units to the desired units. �     	   @ ����       >��>��0�p_?���       	   "DCAT|Control|Waveform Refresh Rate   ms   $Specifies the waveform refresh rate. �            d          DCAT|Data|Async AI Data 1       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 10       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 11       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 12       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 13       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 14       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 15       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 16       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 2       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 3       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 4       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 5       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 6       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 7       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 8       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async AI Data 9       ,Contains the asynchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Async DI Data 1       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 10       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 11       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 12       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 13       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 14       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 15       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 16       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 2       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 3       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 4       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 5       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 6       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 7       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 8       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async DI Data 9       ;Contains the asynchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Async Time 1   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 10   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 11   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 12   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 13   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 14   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 15   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 16   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 2   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 3   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 4   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 5   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 6   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 7   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 8   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Async Time 9   ms   )Contains the asynchronous data timestamp. �     	   @ ����                      	    DCAT|Data|FPGA Data 1       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 10       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 11       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 12       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 13       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 14       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 15       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 16       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 2       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 3       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 4       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 5       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 6       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 7       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 8       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|FPGA Data 9       B"Contains the FPGA ID, Timestamp, and Data the rows of the array." �     	   @ ��������                                 
    DCAT|Data|MS Data 1       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 10       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 11       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 12       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 13       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 14       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 15       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 16       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 2       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 3       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 4       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 5       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 6       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 7       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 8       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Data 9       Contains the medium speed data. �     	   @ ��������                                 
    DCAT|Data|MS Time 1   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 10   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 11   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 12   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 13   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 14   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 15   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 16   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 2   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 3   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 4   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 5   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 6   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 7   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 8   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|MS Time 9   ms   )Contains the medium speed data timestamp. �     	   @ ����                      	    DCAT|Data|Sync AI Data 1       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 10       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 11       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 12       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 13       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 14       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 15       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 16       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 2       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 3       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 4       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 5       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 6       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 7       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 8       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync AI Data 9       +Contains the synchronous analog input data. �     	   @ ��������                                 
    DCAT|Data|Sync DI Data 1       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 10       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 11       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 12       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 13       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 14       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 15       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 16       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 2       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 3       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 4       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 5       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 6       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 7       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 8       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync DI Data 9       :Contains the synchronous digital input data as a bitfield. �     	   @ ����                      	    DCAT|Data|Sync Time 1   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 10   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 11   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 12   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 13   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 14   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 15   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 16   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 2   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 3   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 4   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 5   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 6   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 7   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 8   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    DCAT|Data|Sync Time 9   ms   (Contains the synchronous data timestamp. �     	   @ ����                      	    
DCAT|EPT|A   
True|False   ,Indicates the state of the encoder A signal. �     !               
DCAT|EPT|B   
True|False   ,Indicates the state of the encoder B signal. �     !               DCAT|EPT|Crank Count       IIndicates the current crank count of the engine position tracking system. �                        DCAT|EPT|Crank Count Max       ^Indicates the maximum crank count observed after starting the engine position tracking system. �                        DCAT|EPT|Crank Count Min       ^Indicates the minimum crank count observed after starting the engine position tracking system. �                        DCAT|EPT|Crank Position   CAT   FIndicates the current position of the engine position tracking system. �                        DCAT|EPT|Cycle       OIndicates the current cycle after starting the engine position tracking system. �                        DCAT|EPT|Cycle Period   Ticks   SIndicates the current cycle period measured by the engine position tracking system. �                        DCAT|EPT|FPGA Time   ns   %Indicates the current FPGA timestamp. �                        DCAT|EPT|Gate-Reset   
True|False   5Indicates the state of the encoder Gate/Reset signal. �     !               DCAT|EPT|Max CAT   CAT   OIndicates the maximum crank angle ticks of the engine position tracking system. �                        DCAT|EPT|Overspeed   Overspeed|Speed OK   DIndicates an overspeed state of the engine position tracking system. �     !               DCAT|EPT|Stalled   Stalled|Running   AIndicates a stalled state of the engine position tracking system. �     !               DCAT|EPT|Start Time   ns   ZIndicates the start time of the current DAQ sampling task according to the FPGA timestamp. �                        DCAT|EPT|Sync   Sync|UnSync   FIndicates a synchronized state of the engine position tracking system. �     !               
DCAT|EPT|Z   
True|False   ,Indicates the state of the encoder Z signal. �     !                DCAT|Encoder Debug|Check Encoder   |    Updates the encoder debug scope. �     !              (DCAT|Encoder Debug|Debug Buffer Overflow   |   .Indicates the DCAT Encoder Debug FIFO is full. �     !               %DCAT|Encoder Debug|Encoder Scope Data       9"Z, A, B, and Gate bits along with associated timestamp." �     	   @ ����               	    DCAT|Engine|Actual TDC Offset   CAD   XIndicates the actual top dead center offset used by the engine position tracking system. �     	                   DCAT|Engine|Async Rate   kS/s   3Specifies the sample rate of the asynchronous data. �     	    B�            DCAT|Engine|Bore   m   Specifies the cylinder bore. �     	    =��          DCAT|Engine|Clearance Volume   liter   �Specifies the clearance volume of the cylinder. [Compression Ratio = (Displacement Volume + Clearance Volume) / Clearance Volume] �     	    <�          DCAT|Engine|Compression Ratio       }Indicates the calculated compression ratio. [Compression Ratio = (Displacement Volume + Clearance Volume) / Clearance Volume] �     	    A�             !DCAT|Engine|Connecting Rod Length   m   $Specifies the connecting rod length. �     	    >�          DCAT|Engine|Crown Area   %   ASpecifies the piston crown surface area relative to the bore area �     	    B�            DCAT|Engine|Cycle Resolution   ppc   *Indicates the calculated cycle resolution. �           �           DCAT|Engine|Cylinder Count       .Defines the number of cylinders in the engine. �                      DCAT|Engine|Cylinder TDC   DATDC   UDefines the cylinder Top Dead Center offsets relative to the absolute encoder offset. �     	   @ ����                                                                              	   DCAT|Engine|Digital Filter   us   NDefines the digital glitch filter used by the engine position tracking system. �     	    ?             DCAT|Engine|Displacement Volume   liter   Indicates the calculated displacement volume. [Compression Ratio = (Displacement Volume + Clearance Volume) / Clearance Volume] �     	    >�nN           DCAT|Engine|Dynamic Start-Stop   |   EEnables dynamically starting and stopping the engine while recording. �     !              DCAT|Engine|Encoder Divide       �"Specifies the level to divide the extrapolated resolution by in order to determine the final sample resolution (Not all combinations of encoder resolution, extrapolation level, and encoder divide are valid.)" �                       DCAT|Engine|Encoder Extrap Level       cSpecifies the level of encoder extrapolation used in the engine position tracking system. (2 valid) �                    DCAT|Engine|Encoder Resolution   ppr   OSpecifies the encoder resolution as it is seen by the engine position tracking. �           h          DCAT|Engine|Encoder Setup   'A Rising Edge|A Any Edge|A & B Any Edge   PDetermines which encoder events are used by the engine position tracking system. �                       DCAT|Engine|Encoder Setup Error   Error|   AIndicates an error in the engine position tracking configuration. �     !               DCAT|Engine|Engine       0Specifies the name or description of the engine. �     0����      GM 1.9L Diesel          DCAT|Engine|Exhaust Valve Close   DATDC   2Specifies the nominal exhaust valve closing angle. �     	    C�            DCAT|Engine|Exhaust Valve Open   DATDC   2Specifies the nominal exhaust valve opening angle. �     	    C4            DCAT|Engine|Head Area   %   CSpecifies the cylinder head surface area relative to the bore area. �     	    B�            DCAT|Engine|Intake Valve Close   DATDC   1Specifies the nominal intake valve closing angle. �     	    �4            DCAT|Engine|Intake Valve Open   DATDC   1Specifies the nominal intake valve opening angle. �     	    ô            DCAT|Engine|Max CAT   CAT   PIndicates the maximum crank angle ticks for the engine position tracking system. �           @           DCAT|Engine|Max Speed   RPM   *Specifies the maximum speed of the engine. �     	    E��           DCAT|Engine|Max Sync Rate   kS/s   LSpecifies the maximum sample rate of the synchronous measurement DAQ device. �     	    C�            DCAT|Engine|Medium Speed Rate   S/s   2Specifies the sample rate of the medium speed DAQ. �     	    A             DCAT|Engine|No FPGA   No FPGA (uDCAT)|FPGA (DCAT)   iSpecifies if the system is configured for acquiring data without an FPGA engine position tracking system. �     !              DCAT|Engine|Operator       Specifies the engine operator. �     0����                 DCAT|Engine|Phase   !1 Z/Cycle|Gate Z|Random Z|Reset Z   �Determines the method of preprocessing the encoder signal to pass only a single index pulse per cycle to the engine position tracking system. �                      DCAT|Engine|Pin Offset   m   Specifies the pin offset. �     	                  DCAT|Engine|Polytropic Exponent       >Specifies the nominal polytropic exponent of the cylinder gas. �     	    ?��          &DCAT|Engine|Polytropic Exponent Source   Constant Value|Calculated Value   JSpecifies the source of the polytropic exponent value used in calculations �                       DCAT|Engine|Project       #Specifies the current test project. �     0����                 DCAT|Engine|Random Z   ppr   1Defines which cycle to use when using a random z. �                     $DCAT|Engine|Reduced Cycle Resolution   ppc   2Indicates the calculated reduced cycle resolution. �           �           DCAT|Engine|Reduced Divide       SIndicated the reduced resolution divide required to obtain the reduced resolution.  �                       DCAT|Engine|Reduced Resolution   ppr   ?Indicates the calculated reduced resolution encoder resolution. �           h           DCAT|Engine|Rotations Per Cycle       GDefines the number of rotations per cycle. (2-Stroke = 1; 4-Stroke = 2) �                    DCAT|Engine|Sample Resolution   ppr   IIndicates the calculated sample resolution based on the encoder settings. �           h           DCAT|Engine|Start-Stop Rate   kS/s   dSpecifies the synchronous sample rate while the engine position tracking system is not synchronized. �     	    A             DCAT|Engine|Stroke   m   8Specifies the piston stroke. (Stroke = 2 * Crank Radius) �     	    =�#�          DCAT|Engine|TDC Offset   CAD   �Specifies the global TDC offset. It is commonly used to easily adjust for changes in the encoder without needing to change each cylinder TDC.  �     	                  DCAT|Engine|Volume File Enable   File|Calculations   MEnables use of use of a volume file instead of using the volume calculations. �     !              DCAT|Engine|Volume File Path       =Specifies the volume file to use instead of the calculations. �     0����                 DCAT|Engine|cDAQ DIO Module       LSpecifies the encoder index signal name when using uDCAT and a cDAQ chassis. �     0����                 DCAT|Error|Align Code       #Indicates the Alignment error code. �                        DCAT|Error|Align Error   Error|No Error   Indicates an Alignment error. �     !               DCAT|Error|Align Text       #Indicates the Alignment error text. �     0����                  DCAT|Error|DAQ Code       Indicates the DAQ error code. �                        DCAT|Error|DAQ Error   Error|No Error   Indicates a DAQ error. �     !               DCAT|Error|DAQ Text       Indicates the DAQ error text. �     0����                  DCAT|Error|Display Code       !Indicates the Display error code. �                        DCAT|Error|Display Error   Error|No Error   Indicates a Display error. �     !               DCAT|Error|Display Text       !Indicates the Display error text. �     0����                  DCAT|Error|FPGA Code       Indicates the FPGA error code. �                        DCAT|Error|FPGA Error   Error|No Error   Indicates an FPGA error. �     !               DCAT|Error|FPGA Text       Indicates the FPGA error text. �     0����                  DCAT|Error|Global Error   Error|No Error   Indicates a global error. �     !               DCAT|Error|Next-Cycle Code       $Indicates the Next-Cycle error code. �                        DCAT|Error|Next-Cycle Error   Error|No Error   Indicates a Next-Cycle error. �     !               DCAT|Error|Next-Cycle Text       $Indicates the Next-Cycle error text. �     0����                  DCAT|Error|Process Code       !Indicates the Process error code. �                        DCAT|Error|Process Error   Error|No Error   Indicates a Process error. �     !               DCAT|Error|Process Text       !Indicates the Process error text. �     0����                  DCAT|Error|Raw Code       "Indicates the Raw File error code. �                        DCAT|Error|Raw Error   Error|No Error   Indicates a Raw File error. �     !               DCAT|Error|Raw Text       "Indicates the Raw File error text. �     0����                  DCAT|Error|Summary Code       &Indicates the Summary File error code. �                        DCAT|Error|Summary Error   Error|No Error   Indicates a Summary File error. �     !               DCAT|Error|Summary Text       &Indicates the Summary File error text. �     0����                  DCAT|Execution|Basic   us   )Execution time of the Basic calculations. �                        DCAT|Execution|Calibrate   us   -Execution time of the Calibrate calculations. �                        DCAT|Execution|Cam   us   'Execution time of the Cam calculations. �                        DCAT|Execution|FPGA   us   (Execution time of the FPGA calculations. �                        DCAT|Execution|Filter   us   *Execution time of the Filter calculations. �                        DCAT|Execution|Gas Temp   us   3Execution time of the Gas Temperature calculations. �                        DCAT|Execution|Heat Release   us   0Execution time of the Heat Release calculations. �                        DCAT|Execution|Injector   us   ,Execution time of the Injector calculations. �                        DCAT|Execution|Knock   us   )Execution time of the Knock calculations. �                        DCAT|Execution|MEP   us   ;Execution time of the Mean Effective Pressure calculations. �                        DCAT|Execution|Medium Speed   us   0Execution time of the Medium Speed calculations. �                        DCAT|Execution|Misfire   us   +Execution time of the Misfire calculations. �                        DCAT|Execution|Motoring   us   ,Execution time of the Motoring calculations. �                        DCAT|Execution|Noise   us   )Execution time of the Noise calculations. �                        DCAT|Execution|PWM   us   :Execution time of the Pulse Width Modulation calculations. �                        DCAT|Execution|Pegging   us   +Execution time of the Pegging calculations. �                        DCAT|Execution|Pump   us   4Execution time of the Synchronous Pump calculations. �                        DCAT|Execution|Scale   us   &Execution time of the Scaling process. �                        DCAT|Execution|Separate   us   )Execution time of the Separating process. �                        DCAT|Execution|Spark   us   )Execution time of the Spark calculations. �                        DCAT|Execution|TDC Offset   us   1Execution time of the TDC Offset Fine Adjustment. �                         DCAT|Execution|User Calculations   us   (Execution time of the User calculations. �                        DCAT|Execution|User Process   us   #Execution time of the User process. �                        DCAT|FPGA|Gain       &Gain associated with each measurement. �     	   @ ����               	   DCAT|FPGA|ID       )ID associated with each FPGA measurement. �     	   @ ����               	   DCAT|FPGA|Name       5Name or description associated with each measurement. �     0����                 DCAT|FPGA|Offset       (Offset associated with each measurement. �     	   @ ����               	   DCAT|FPGA|Units       'Units associated with each measurement. �     0����                 DCAT|Filter|Filter        Defines the type of filter used. �     	   @ ����                                                                              	   DCAT|Filter|Frequency   %   |Defines the filter frequency as a percent of the nyquist frequency. This value is only valid when using FIR and IIR filters. �     	   @ ����                                                                              	   DCAT|Filter|N       yDefines the number of cycles to include in the rolling average or the number of samples to include in the boxcar average. �     	   @ ����                                                                              	   DCAT|Filter|Order       CDefines the order of the filter when using the FIR and IIR filters. �     	   @ ����                                                                              	   DCAT|HR|C1c       8Woschni Coefficient 1 for Compression  (Default = 2.28). �     	    @�          DCAT|HR|C1e       DWoschni Coefficient 1 for Combustion and Expansion (Default = 2.28). �     	    @�          DCAT|HR|C1ge       8Woschni Coefficient 1 for Gas Exchange (Default = 6.18). �     	    @�          DCAT|HR|C2c       6Woschni Coefficient 2 for Compression (Default = 0.0). �     	                  DCAT|HR|C2e       GWoschni Coefficient 2 for Combustion and Expansion (Default = 0.00324). �     	    ;TV.          DCAT|HR|C2ge       7Woschni Coefficient 2 for Gas Exchange (Default = 0.0). �     	                  DCAT|HR|End Angle   CAD   <Specifies the angle to end looking for the end of combustion �     	    Bp            DCAT|HR|End of Combustion   /Constant|N Below Zero|Boxcar Average Below Zero   =Specifies the method used to determine the end of combustion. �                       DCAT|HR|Heat Release   �Single Zone|Single Zone Dual Transducer|Single Zone + Heat Transfer|Single Zone Dual Transducer + Heat Transfer|Modified Rassweiler and Withrow|Pressure Ratio|User Defined   4Specifies the method used to calculate heat release. �                       DCAT|HR|Heat Transfer   W/m2-K   SDefines the heat transfer when using the constant Heat Transfer Correlation method. �     	                  !DCAT|HR|Heat Transfer Correlation   ,Constant|Woschni 1978|Woschni 1990|Hohenberg   ESpecifies the method used to calculate the Heat Transfer Correlation. �                       DCAT|HR|N End       NSpecifies the number of samples to use when determining the end of combustion. �                      DCAT|HR|N Start       PSpecifies the number of samples to use when determining the start of combustion. �                      DCAT|HR|Polytropic Correlation   LHayes (SAE860029)|Indolene (SAE841359)|Propane (SAE841359)|Custom (a*T(K)+b)   >Specifies the method use to calculate the polytropic exponent. �                       DCAT|HR|PreChamber Volume   liter   LSpecifies the volume of the prechamber used in dual transducer calculations. �     	                  DCAT|HR|Smoothing   %   DPressure waveform smoothing factor as a percent of one engine cycle. �     	    ?�            DCAT|HR|Start Angle   CAD   @Specifies the angle to start looking for the start of combustion �     	    ��            DCAT|HR|Start of Combustion   VConstant|N Below Zero|Boxcar Average Below Zero|N Above Zero|Boxcar Average Above Zero   ?Specifies the method used to determine the start of combustion. �                       DCAT|HR|Wall Temperature   K   PSpecifies the Wall Temperature when using the constant Wall Temperature Profile. �     	    C��           DCAT|HR|Wall Temperature BDC   K   aSpecifies the Bottom Dead Center Wall Temperature when using the linear Wall Temperature Profile. �     	    C��            DCAT|HR|Wall Temperature Profile   Constant|Linear   MSpecifies the method used to calculate the cylinder Wall Temperature Profile. �                       DCAT|HR|Wall Temperature TDC   K   ^Specifies the Top Dead Center Wall Temperature when using the linear Wall Temperature Profile. �     	    C��           	DCAT|HR|a       c"Defines the Polytropic Exponent Correlation ""a"" Value when using custom Polytropic Correlation." �     	                  	DCAT|HR|b   liter   c"Defines the Polytropic Exponent Correlation ""b"" Value when using custom Polytropic Correlation." �     	                  !DCAT|Injection|Fuel Rail Pressure   CAD   0Defines the fuel rail pressure of the injectors. �     	                  (DCAT|Injection|Fuel Rail Pressure Source   Constant Value|DAQ Channel   NDetermines the source of the fuel rail pressure used in determining fuel flow. �                       DCAT|Injection|Min Injection   ms   $Defines the minimum injection width. �     	    =���          DCAT|Injection|Signal   Voltage|Current   !Defines the injector signal type. �                       DCAT|Injection|Type   PFI|DI Solenoid|DI Piezo   Defines the injector type. �                       DCAT|Injection|X-Fuel Pressure   MPa   HDefines the X-Axis (Fuel Pressure) of the 2d injector calibration table. �     	   @ ����           ?�         	   DCAT|Injection|Y-Duration   ms   CDefines the Y-Axis (Duration) of the 2d injector calibration table. �     	   @ ����           ?�         	   DCAT|Injection|Z-Fuel Flow   mg/Inj   DDefines the Z-Axis (Fuel Flow) of the 2d injector calibration table. �     	   @ ��������                                 
    DCAT|Knock|High Cutoff Frequency   kHz   JSpecifies the High Cutoff Frequency of the knock filter for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Knock End   CAD   DSpecifies the crank angle to end the knock window for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Knock Start   CAD   FSpecifies the crank angle to start the knock window for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Low Cutoff Frequency   kHz   ISpecifies the Low Cutoff Frequency of the knock filter for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Minimum Reference       MSpecifies the Minimum Reference Value used to remove noise for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Reference End   CAD   HSpecifies the crank angle to end the reference window for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Reference Start   CAD   JSpecifies the crank angle to start the reference window for each cylinder. �     	   @ ����                                                                              	   DCAT|Knock|Threshold       0Specifies the knock threshold for each cylinder. �     	   @ ����                                                                              	   DCAT|Loop|Align Count       4Indicate the current cycles count of the Align loop. �                        DCAT|Loop|Align Period   ms   2Indicate the approximate Period of the Align loop. �     	                   DCAT|Loop|Align Time   ms   2Indicate the time used to complete the Align loop. �     	                   DCAT|Loop|DAQ Count       2Indicate the current cycles count of the DAQ loop. �                        DCAT|Loop|DAQ Period   ms   0Indicate the approximate Period of the DAQ loop. �     	                   DCAT|Loop|DAQ Time   ms   0Indicate the time used to complete the DAQ loop. �     	                   DCAT|Loop|Display Count       6Indicate the current cycles count of the Display loop. �                        DCAT|Loop|Display Period   ms   4Indicate the approximate Period of the Display loop. �     	                   DCAT|Loop|Display Time   ms   4Indicate the time used to complete the Display loop. �     	                   DCAT|Loop|FPGA Control Count       ;Indicate the current cycles count of the FPGA Control loop. �                        DCAT|Loop|FPGA Control Period   ms   9Indicate the approximate Period of the FPGA Control loop. �     	                   DCAT|Loop|FPGA Control Time   ms   9Indicate the time used to complete the FPGA Control loop. �     	                   "DCAT|Loop|Next-Cycle Control Count       AIndicate the current cycles count of the Next-Cycle Control loop. �                        #DCAT|Loop|Next-Cycle Control Period   ms   ?Indicate the approximate Period of the Next-Cycle Control loop. �     	                   !DCAT|Loop|Next-Cycle Control Time   ms   ?Indicate the time used to complete the Next-Cycle Control loop. �     	                   DCAT|Loop|Process Count       6Indicate the current cycles count of the Process loop. �                        DCAT|Loop|Process Period   ms   4Indicate the approximate Period of the Process loop. �     	                   DCAT|Loop|Process Time   ms   4Indicate the time used to complete the Process loop. �     	                   DCAT|Loop|Raw File Count       7Indicate the current cycles count of the Raw File loop. �                        DCAT|Loop|Raw File Period   ms   5Indicate the approximate Period of the Raw File loop. �     	                   DCAT|Loop|Raw File Time   ms   5Indicate the time used to complete the Raw File loop. �     	                   DCAT|Loop|Summary File Count       ;Indicate the current cycles count of the Summary File loop. �                        DCAT|Loop|Summary File Period   ms   9Indicate the approximate Period of the Summary File loop. �     	                   DCAT|Loop|Summary File Time   ms   9Indicate the time used to complete the Summary File loop. �     	                   DCAT|Medium Speed|CJC Channel       {Cold junction compensation channel associated with each measurement when using a channel cold junction compensation source. �     0����                 DCAT|Medium Speed|CJC Source       CCold junction compensation source associated with each measurement. �     	   @ ����               	   DCAT|Medium Speed|CJC Value       zCold junction compensation value associated with each measurement when using a constant cold junction compensation source. �     	   @ ����               	   DCAT|Medium Speed|Disable       LDisables data acquisition and calculations associated with each measurement. �     	   @ ����               	   DCAT|Medium Speed|Filter Cutoff       !Knock Threshold for Each Cylinder �     	   @ ����               	   DCAT|Medium Speed|Gain       &Gain associated with each measurement. �     	   @ ����               	   DCAT|Medium Speed|Max       L"Maximum voltage, current, or temperature associated with each measurement." �     	   @ ����               	   DCAT|Medium Speed|Min       L"Minimum voltage, current, or temperature associated with each measurement." �     	   @ ����               	   DCAT|Medium Speed|Name       5Name or description associated with each measurement. �     0����                 DCAT|Medium Speed|Offset       (Offset associated with each measurement. �     	   @ ����               	   "DCAT|Medium Speed|Physical Channel       2Physical channel associated with each measurement. �     0����                 DCAT|Medium Speed|Save Trigger       sEnables the channel to be used to trigger the start of a file save. Each index is associated with each measurement. �     	   @ ����               	   DCAT|Medium Speed|Scaling       0Scaling method associated with each measurement. �     	   @ ����               	   (DCAT|Medium Speed|Terminal Configuration       8Terminal configuration associated with each measurement. �     	   @ ����               	   #DCAT|Medium Speed|Thermocouple Type       3Thermocouple type associated with each measurement. �     	   @ ����               	   DCAT|Medium Speed|Units       'Units associated with each measurement. �     0����                 DCAT|Misfire|Misfire   =Peak Pressure|Net Mean Effective Pressure|Combustion Pressure   2Specifies the method to use for Misfire detection. �                       DCAT|Misfire|Threshold   kPa   jSpecifies the threshold used to detect a misfire. The use of the value depends on the misfire method used. �     	    Dz            DCAT|Next-Cycle|Basic   Enabled|Disabled   6Enables the Basic calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Cam   Enabled|Disabled   4Enables the Cam calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|FPGA   Enabled|Disabled   5Enables the FPGA calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Gas Temp   Enabled|Disabled   @Enables the Gas Temperature calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Heat Release   Enabled|Disabled   =Enables the Heat Release calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Injector   Enabled|Disabled   9Enables the Injector calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Knock   Enabled|Disabled   6Enables the Knock calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|MEP   Enabled|Disabled   HEnables the Mean Effective Pressure calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Medium Speed   Enabled|Disabled   =Enables the Medium Speed calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Misfire   Enabled|Disabled   8Enables the Misfire calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Motoring   Enabled|Disabled   9Enables the Motoring calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Noise   Enabled|Disabled   6Enables the Noise calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|PWM   Enabled|Disabled   GEnables the Pulse Width Modulation calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Pump   Enabled|Disabled   AEnables the Synchronous Pump calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|Spark   Enabled|Disabled   6Enables the Spark calculations for Next-Cycle control. �     !             !DCAT|Next-Cycle|User Calculations   Enabled|Disabled   5Enables the User calculations for Next-Cycle control. �     !             DCAT|Next-Cycle|User Process   Enabled|Disabled   3Enables the User Processing for Next-Cycle control. �     !              DCAT|Pegging|Location   CAD   eSpecifies the location used to peg cylinder pressure when using constant and synchronous MAP pegging. �     	    Ö            DCAT|Pegging|Pegging   (None|Constant|Synchronous MAP|Polytropic   3Specifies the method used to peg cylinder pressure. �                       DCAT|Pegging|Pegging Pressure   kPa abs   QSpecifies the pressure used to peg cylinder pressure when using constant pegging. �     	    B�             DCAT|Pegging|Polytropic Exponent       >Specifies the polytropic exponent used for polytropic pegging. �     	    ?��          DCAT|Pegging|Window   CAD   WThe crank angle window size used to average noise in synchronous waveform measurements. �     	    @�            DCAT|Raw|Comments       +User comments to be included in data files. �     0����                 DCAT|Raw|Continuous   Continuous|Single   rDetermines if the logging process will stop after a single point or automatically start a new point when finished. �     !              DCAT|Raw|Cycle Limit       9Specifies the maximum cycle count of a file when enabled. �                       DCAT|Raw|Enable Cycle Limit   Cycle Limit|No Cycle Limit   )Enables the cycle limit for file logging. �     !              DCAT|Raw|Enable Size Limit   Size Limit|No Size Limit   (Enables the size limit for file logging. �     !              DCAT|Raw|Enable Time Limit   Time Limit|No Time Limit   (Enables the time limit for file logging. �     !              DCAT|Raw|Error   Error|No Error   (Indicates a Raw File post process error. �     !               DCAT|Raw|Error Code       /Indicates the Raw File post process error code. �                        DCAT|Raw|Error Text       2Indicates the Raw File post processing error text. �     0����                  DCAT|Raw|File       !Current raw data file processing. �     0����                  DCAT|Raw|File Counter       -Indicates the file count of the current file. �                        DCAT|Raw|File Name       j"Raw file name. Use general time format to insert a timestamp. Use ""XXX"" to insert file counter number." �     0����      Raw_XXX          DCAT|Raw|File Part       2Indicates the part of the current continuous file. �                        DCAT|Raw|File Path       .Indicates the path of the current saving file. �     0����                  DCAT|Raw|File Progress   %   +Indicates the progress of the current file. �     	                   DCAT|Raw|Overwrite File   Overwrite|New File   JIndicates if a file will be overwritten during the next file save process. �     !               DCAT|Raw|Path       )Specifies the folder for saving raw data. �     0����      C:\Data          DCAT|Raw|Process File       $Defines the summary post process VI. �     0����                 DCAT|Raw|Queue       7Array of file names in the Raw File post process queue. �     0����                  DCAT|Raw|Reset Counter   Reset Counter|   3Resets the file counter to a user specified number. �     !              DCAT|Raw|Reset Counter Value        Value to reset the file counter. �                       DCAT|Raw|Save Trigger   MS Save Trigger|Manual Trigger   EEnables starting file saving events from a medium speed save trigger. �     !              DCAT|Raw|Saving File   Saving|Standby   AIndicates that a file is currently in the process of being saved. �     !               DCAT|Raw|Size Limit   MB   2Specifies the maximum size of a file when enabled. �     	                  DCAT|Raw|Start-Stop File   Start or Stop File|   'Starts or stops a file logging process. �     !              DCAT|Raw|Time Limit   s   9Specifies the maximum record time of a file when enabled. �     	                  DCAT|Results|Avaliable Results       ?Indicates the available statistical results calculated by DCAT. �     0����                  DCAT|Results|Cycle       "Indicates the current cycle count. �                        DCAT|Results|Speed   RPM   #Indicates the current engine speed. �     	                   DCAT|Results|Time   ns   2Indicates the current timestamp of the FPGA timer. �                        DCAT|Separate|Conversion   Fast|Accurate   KSpecifies the method used to convert synchronous data to asynchronous data. �                       DCAT|Simulation|Cam Duration   CAD   %Specifies the simulated cam duration. �     	   @ ����       BH  C>  C>         	   DCAT|Simulation|Cam Start   CAD   "Specifies the simulated cam start. �     	   @ ����       �  B�  C�         	   DCAT|Simulation|Exhaust Cam   CAD   +Specifies the simulated exhaust cam offset. �     	                  "DCAT|Simulation|Fuel Rail Pressure   MPa abs   +Specifies the simulated fuel rail pressure. �     	    A             "DCAT|Simulation|Injection Duration   ms   +Specifies the simulated injection duration. �     	   @ ����       >���?���       	   "DCAT|Simulation|Injection Location   CAD   +Specifies the simulated injection locations �     	   @ ����       ��  �          	   DCAT|Simulation|Intake Cam   CAD   *Specifies the simulated intake cam offset. �     	                  *DCAT|Simulation|Manifold Absolute Pressure   kPa abs   3Specifies the simulated manifold absolute pressure. �     	    B�            DCAT|Simulation|PWM Duty Cycle   %   <Specifies the simulated pulse width  measurement duty cycle. �     	    BH            DCAT|Simulation|PWM Frequency   kHz   ;Specifies the simulated pulse width  measurement frequency. �     	    A             DCAT|Simulation|Spark Dwell   ms   $Specifies the simulated spark dwell. �     	    ?�            DCAT|Simulation|Spark Location   CAD   'Specifies the simulated spark location. �     	   @ ����       ¾  ��         	   DCAT|Simulation|Speed   RPM   %Specifies the simulated engine speed. �     	    Dz            )DCAT|Simulation|Synchronous Pump Duration   CAD   2Specifies the simulated synchronous pump duration. �     	    BH            &DCAT|Simulation|Synchronous Pump Start   CAD   /Specifies the simulated synchronous pump start. �     	   @ ����       Ö  �p  C4         	   DCAT|Spark|Min Dwell   ms    Defines the minimum dwell width. �     	    =���          DCAT|Spark|Restrike Delay   ms   #Defines the maximum restrike delay. �     	    ?�            DCAT|Spark|Signal   Voltage|Current   Defines the spark signal type. �                       #DCAT|Statistics|Basic Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    #DCAT|Statistics|Basic Results Names       *Contains the names of the rolling results. �     0����                  !DCAT|Statistics|Cam Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    !DCAT|Statistics|Cam Results Names       *Contains the names of the rolling results. �     0����                  #DCAT|Statistics|Cycle Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    #DCAT|Statistics|Cycle Results Names       *Contains the names of the rolling results. �     0����                  "DCAT|Statistics|FPGA Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    "DCAT|Statistics|FPGA Results Names       *Contains the names of the rolling results. �     0����                  *DCAT|Statistics|Heat Release Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    *DCAT|Statistics|Heat Release Results Names       *Contains the names of the rolling results. �     0����                  'DCAT|Statistics|Injection Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    'DCAT|Statistics|Injection Results Names       *Contains the names of the rolling results. �     0����                  #DCAT|Statistics|Knock Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    #DCAT|Statistics|Knock Results Names       *Contains the names of the rolling results. �     0����                  !DCAT|Statistics|MEP Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    !DCAT|Statistics|MEP Results Names       *Contains the names of the rolling results. �     0����                  *DCAT|Statistics|Medium Speed Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    *DCAT|Statistics|Medium Speed Results Names       *Contains the names of the rolling results. �     0����                  %DCAT|Statistics|Misfire Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    %DCAT|Statistics|Misfire Results Names       *Contains the names of the rolling results. �     0����                  #DCAT|Statistics|Noise Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    #DCAT|Statistics|Noise Results Names       *Contains the names of the rolling results. �     0����                  !DCAT|Statistics|PWM Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    !DCAT|Statistics|PWM Results Names       *Contains the names of the rolling results. �     0����                  %DCAT|Statistics|Pegging Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    %DCAT|Statistics|Pegging Results Names       *Contains the names of the rolling results. �     0����                  "DCAT|Statistics|Pump Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    "DCAT|Statistics|Pump Results Names       *Contains the names of the rolling results. �     0����                  (DCAT|Statistics|Slow Speed Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    (DCAT|Statistics|Slow Speed Results Names       *Contains the names of the rolling results. �     0����                  #DCAT|Statistics|Spark Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    #DCAT|Statistics|Spark Results Names       *Contains the names of the rolling results. �     0����                  "DCAT|Statistics|User Results Array       WContains the results of the calculations and rolling statistics for those calculations. �     	   @ ��������                                 
    "DCAT|Statistics|User Results Names       *Contains the names of the rolling results. �     0����                  DCAT|Sum|Comments       +User comments to be included in data files. �     0����                 DCAT|Sum|Continuous   Continuous|Single   rDetermines if the logging process will stop after a single point or automatically start a new point when finished. �     !              DCAT|Sum|Cycle Limit       9Specifies the maximum cycle count of a file when enabled. �                       DCAT|Sum|Enable Cycle Limit   Cycle Limit|No Cycle Limit   )Enables the cycle limit for file logging. �     !              DCAT|Sum|Enable Size Limit   Size Limit|No Size Limit   (Enables the size limit for file logging. �     !              DCAT|Sum|Enable Time Limit   Time Limit|No Time Limit   (Enables the time limit for file logging. �     !              DCAT|Sum|Error   Error|No Error   /Indicates a Summary File post processing error. �     !               DCAT|Sum|Error Code       6Indicates the Summary File post processing error code. �                        DCAT|Sum|Error Text       3Indicates the Summary File post process error text. �     0����                  DCAT|Sum|File       %Current summary data file processing. �     0����                  DCAT|Sum|File Counter       -Indicates the file count of the current file. �                        DCAT|Sum|File Name       n"Summary file name. Use general time format to insert a timestamp. Use ""XXX"" to insert file counter number." �     0����      Sum_XXX          DCAT|Sum|File Part       2Indicates the part of the current continuous file. �                        DCAT|Sum|File Path       .Indicates the path of the current saving file. �     0����                  DCAT|Sum|File Progress   %   +Indicates the progress of the current file. �     	                   DCAT|Sum|Overwrite File   Overwrite|New File   JIndicates if a file will be overwritten during the next file save process. �     !               DCAT|Sum|Path       -Specifies the folder for saving summary data. �     0����      C:\Data          DCAT|Sum|Process File       $Defines the summary post process VI. �     0����                 DCAT|Sum|Queue       ;Array of file names in the Summary File post process queue. �     0����                  DCAT|Sum|Reset Counter   Reset Counter|   3Resets the file counter to a user specified number. �     !              DCAT|Sum|Reset Counter Value        Value to reset the file counter. �                       DCAT|Sum|Save Trigger   MS Save Trigger|Manual Trigger   EEnables starting file saving events from a medium speed save trigger. �     !              DCAT|Sum|Saving File   Saving|Standby   AIndicates that a file is currently in the process of being saved. �     !               DCAT|Sum|Size Limit   MB   2Specifies the maximum size of a file when enabled. �     	                  DCAT|Sum|Start-Stop File   Start or Stop File|   'Starts or stops a file logging process. �     !              DCAT|Sum|Time Limit   s   9Specifies the maximum record time of a file when enabled. �     	                  DCAT|Sync Digital|Cylinder       9Cylinders associated with each measurement in a bitfield. �     	   @ ����       G� G� G� G�                                                        	   DCAT|Sync Digital|Invert       <Invert the digital signals associated with each measurement. �     	   @ ����                                                                              	   DCAT|Sync Digital|Name       &Name associated with each measurement. �     0����      gTDC;Data;Reduce Resolution;Reserved;DI 4;DI 5;DI 6;DI 7;DI 8;DI 9;DI 10;DI 11;DI 12;DI 13;DI 14;DI 15
          DCAT|Sync Digital|Type       2Measurement Type associated with each measurement. �     	   @ ����                                                                              	   DCAT|Sync|Cylinder       9Cylinders associated with each measurement in a bitfield. �     	   @ ����               	   DCAT|Sync|Disable       LDisables data acquisition and calculations associated with each measurement. �     	   @ ����               	   DCAT|Sync|Filter       HFilter resource number associated with each measurement. (0 = No Filter) �     	   @ ����               	   DCAT|Sync|Gain       cGain associated with each measurement when using  the gain only or gain and offset scaling methods. �     	   @ ����               	   DCAT|Sync|Max       ?Maximum channel voltage range associated with each measurement. �     	   @ ����               	   DCAT|Sync|Min       ?Minimum channel voltage range associated with each measurement. �     	   @ ����               	   DCAT|Sync|Name       5Name or description associated with each measurement. �     0����                 DCAT|Sync|Offset       VOffset associated with each measurement when using the gain and offset scaling method. �     	   @ ����               	   DCAT|Sync|Physical Channel       2Physical channel associated with each measurement. �     0����                 !DCAT|Sync|Polynomial Coefficients       bPolynomial Coefficients associated with each measurement when using the polynomial scaling method. �     	   @ ��������                         
   DCAT|Sync|Scaling       0Scaling method associated with each measurement. �     	   @ ����               	   DCAT|Sync|Table X       STable X array associated with each measurement when using the table scaling method. �     	   @ ��������                         
   DCAT|Sync|Table Y       STable Y array associated with each measurement when using the table scaling method. �     	   @ ��������                         
    DCAT|Sync|Terminal Configuration       >Terminal Configuration array associated with each measurement. �     	   @ ����               	   DCAT|Sync|Type       2Measurement Type associated with each measurement. �     	   @ ����               	   DCAT|Sync|Units       'Units associated with each measurement. �     0����                 DCAT|System|CPU   %   >Indicates the average CPU use of the system. (RT Systems Only) �     	    B��           DCAT|System|Core   %   LIndicates the current CPU use for each core in the system. (RT Systems Only) �     	   @ ����       B���B�2�       	    DCAT|System|DAQmx       `This array represents the DAQmx configuration of the system flattened to an array of characters. �     	   @ ����      �      Dev1�lf  94  1'   PXI-6123          Dev1/ai0   Dev1/ai1   Dev1/ai2   Dev1/ai3   Dev1/ai4   Dev1/ai5   Dev1/ai6   Dev1/ai7   
  '�  (&  (<  (=  (>  (?  (R  (S  9�  >lA��    A��       ��      ?�      �      @      �      @      �$      @$                Dev1/port0/line0   Dev1/port0/line1   Dev1/port0/line2   Dev1/port0/line3   Dev1/port0/line4   Dev1/port0/line5   Dev1/port0/line6   Dev1/port0/line7                      Dev1/port0/line0   Dev1/port0/line1   Dev1/port0/line2   Dev1/port0/line3   Dev1/port0/line4   Dev1/port0/line5   Dev1/port0/line6   Dev1/port0/line7   Dev2�le  94  1'   PXI-6123          Dev2/ai0   Dev2/ai1   Dev2/ai2   Dev2/ai3   Dev2/ai4   Dev2/ai5   Dev2/ai6   Dev2/ai7   
  '�  (&  (<  (=  (>  (?  (R  (S  9�  >lA��    A��       ��      ?�      �      @      �      @      �$      @$                Dev2/port0/line0   Dev2/port0/line1   Dev2/port0/line2   Dev2/port0/line3   Dev2/port0/line4   Dev2/port0/line5   Dev2/port0/line6   Dev2/port0/line7                      Dev2/port0/line0   Dev2/port0/line1   Dev2/port0/line2   Dev2/port0/line3   Dev2/port0/line4   Dev2/port0/line5   Dev2/port0/line6   Dev2/port0/line7   Dev3kV  93  1'   PXI-6251          Dev3/ai0   Dev3/ai1   Dev3/ai2   Dev3/ai3   Dev3/ai4   Dev3/ai5   Dev3/ai6   Dev3/ai7   Dev3/ai8   Dev3/ai9   	Dev3/ai10   	Dev3/ai11   	Dev3/ai12   	Dev3/ai13   	Dev3/ai14   	Dev3/ai15   
  '�  (&  (<  (=  (>  (?  (G  (R  (S  >l A3�    A.��       ��������?��������ə�����?ə�������      ?�      ��      ?�      �       @       �      @      �$      @$                Dev3/port0/line0   Dev3/port0/line1   Dev3/port0/line2   Dev3/port0/line3   Dev3/port0/line4   Dev3/port0/line5   Dev3/port0/line6   Dev3/port0/line7   Dev3/port1/line0   Dev3/port1/line1   Dev3/port1/line2   Dev3/port1/line3   Dev3/port1/line4   Dev3/port1/line5   Dev3/port1/line6   Dev3/port1/line7   Dev3/port2/line0   Dev3/port2/line1   Dev3/port2/line2   Dev3/port2/line3   Dev3/port2/line4   Dev3/port2/line5   Dev3/port2/line6   Dev3/port2/line7      Dev3/ao0   Dev3/ao1     (R   �      @      �$      @$                Dev3/port0/line0   Dev3/port0/line1   Dev3/port0/line2   Dev3/port0/line3   Dev3/port0/line4   Dev3/port0/line5   Dev3/port0/line6   Dev3/port0/line7   Dev3/port1/line0   Dev3/port1/line1   Dev3/port1/line2   Dev3/port1/line3   Dev3/port1/line4   Dev3/port1/line5   Dev3/port1/line6   Dev3/port1/line7   Dev3/port2/line0   Dev3/port2/line1   Dev3/port2/line2   Dev3/port2/line3   Dev3/port2/line4   Dev3/port2/line5   Dev3/port2/line6   Dev3/port2/line7   SC1Mod1      9D  1(   	SCXI-1102           SC1Mod1/ai0   SC1Mod1/ai1   SC1Mod1/ai2   SC1Mod1/ai3   SC1Mod1/ai4   SC1Mod1/ai5   SC1Mod1/ai6   SC1Mod1/ai7   SC1Mod1/ai8   SC1Mod1/ai9   SC1Mod1/ai10   SC1Mod1/ai11   SC1Mod1/ai12   SC1Mod1/ai13   SC1Mod1/ai14   SC1Mod1/ai15   SC1Mod1/ai16   SC1Mod1/ai17   SC1Mod1/ai18   SC1Mod1/ai19   SC1Mod1/ai20   SC1Mod1/ai21   SC1Mod1/ai22   SC1Mod1/ai23   SC1Mod1/ai24   SC1Mod1/ai25   SC1Mod1/ai26   SC1Mod1/ai27   SC1Mod1/ai28   SC1Mod1/ai29   SC1Mod1/ai30   SC1Mod1/ai31   	  '�  (&  (<  (=  (>  (?  (R  (S  >l                    ��������?��������$      @$                                     SC1Mod2      9D  1(   
SCXI-1102B           SC1Mod2/ai0   SC1Mod2/ai1   SC1Mod2/ai2   SC1Mod2/ai3   SC1Mod2/ai4   SC1Mod2/ai5   SC1Mod2/ai6   SC1Mod2/ai7   SC1Mod2/ai8   SC1Mod2/ai9   SC1Mod2/ai10   SC1Mod2/ai11   SC1Mod2/ai12   SC1Mod2/ai13   SC1Mod2/ai14   SC1Mod2/ai15   SC1Mod2/ai16   SC1Mod2/ai17   SC1Mod2/ai18   SC1Mod2/ai19   SC1Mod2/ai20   SC1Mod2/ai21   SC1Mod2/ai22   SC1Mod2/ai23   SC1Mod2/ai24   SC1Mod2/ai25   SC1Mod2/ai26   SC1Mod2/ai27   SC1Mod2/ai28   SC1Mod2/ai29   SC1Mod2/ai30   SC1Mod2/ai31   	  '�  (&  (<  (=  (>  (?  (R  (S  >l                    ��������?��������$      @$                                             	    DCAT|System|DCAT License   +Unlicensed|Evaluation|Processing|uDCAT|DCAT   (Indicates the state of the DCAT License. �                        DCAT|System|DCAT Version       Indicates the DCAT version. �     0����      3.120.11300           DCAT|System|Free Disk Space   MB   2Indicates the total free disk space of the system. �     	    Hh��           DCAT|System|RAM   MB   <Indicates the available RAM of the system. (RT Systems Only) �     	    D�p�           DCAT|TDC Offset|Loss Angle   CAD   �Specifies the difference between peak cylinder pressure and cylinder TDC due to heat transfer losses; commonly referred to as the thermodynamic loss angle. �     	    ?             DCAT|TDC Offset|PolyC High       @Sets the upper limit for the polytropic compression coefficient. �     	    ?�=q          DCAT|TDC Offset|PolyC Low       @Sets the lower limit for the polytropic compression coefficient. �     	    ?��          DCAT|TDC Offset|PolyE High       >Sets the upper limit for the polytropic expansion coefficient. �     	    ?�33          DCAT|TDC Offset|PolyE Low       >Sets the lower limit for the polytropic expansion coefficient. �     	    ?�ff          "DCAT|TDC Offset|Reference Cylinder       :Specifies the cylinder used as a reference for TDC offset. �     	    ?�            DCAT|TDC Offset|TDC Fine Adjust   CAD   \Specifies the TDC fine adjustment. A TDC offset may force resampling data which can be slow. �     	                  DCAT|TDC Offset|dPoly High       bSets the upper limit for the difference between polytropic compression and expansion coefficients. �     	    ?             DCAT|TDC Offset|dPoly Low       bSets the lower limit for the difference between polytropic compression and expansion coefficients. �     	    �             DCAT|Temp|Exhaust Pressure   kPa abs   /Pressure of the intake gas at the intake valve. �     	    B�            DCAT|Temp|Exhaust Temperature   K   4Temperature of the exhaust gas at the exhaust valve. �     	    C�            DCAT|Temp|Intake Pressure   kPa abs   1Pressure of the exhaust gas at the exhaust valve. �     	    B�            DCAT|Temp|Intake Temperature   K   2Temperature of the intake gas at the intake valve. �     	    C�            DCAT|Temp|Residual Fraction   Fraction   TFraction of exhaust gas remaining in the combustion chamber after the exhaust event. �     	                  DCAT|Temp|Window   CAD   WThe crank angle window size used to average noise in synchronous waveform measurements. �     	    @�            DCAT|User|User Calculation VI       "Specifies the user calculation VI. �     0����                 DCAT|User|User Heat Release VI       #Specifies the user heat release VI. �     0����                 DCAT|User|User Process VI       !Specifies the user processing VI. �     0����                 DCAT|Waveforms|Acoustic       vWaveform array representing the acoustic signal at each point in the asynchronous sample resolution for each cylinder. �     	   @ ��������                     
    $DCAT|Waveforms|Async Encoder Indexes       vWaveform array representing the asynchronous indexes at each point in the reduced sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Crank Angle   CAD   SWaveform array representing the crank angle at each point in the sample resolution. �     	   @ ����      �ô  ó� ó  ò� ò  ñ� ñ  ð� ð  ï� ï  î� î  í� í  ì� ì  ë� ë  ê� ê  é� é  è� è  ç� ç  æ� æ  å� å  ä� ä  ã� ã  â� â  á� á  à� à  ß� ß  Þ� Þ  Ý� Ý  Ü� Ü  Û� Û  Ú� Ú  Ù� Ù  Ø� Ø  ×� ×  Ö� Ö  Õ� Õ  Ô� Ô  Ó� Ó  Ò� Ò  Ñ� Ñ  Ð� Ð  Ï� Ï  Î� Î  Í� Í  Ì� Ì  Ë� Ë  Ê� Ê  É� É  È� È  Ç� Ç  Æ� Æ  Å� Å  Ä� Ä  Ã� Ã  Â� Â  Á� Á  À� À  �  �~  �}  �|  �{  �z  �y  �x  �w  �v  �u  �t  �s  �r  �q  �p  �o  �n  �m  �l  �k  �j  �i  �h  �g  �f  �e  �d  �c  �b  �a  �`  �_  �^  �]  �\  �[  �Z  �Y  �X  �W  �V  �U  �T  �S  �R  �Q  �P  �O  �N  �M  �L  �K  �J  �I  �H  �G  �F  �E  �D  �C  �B  �A  �@  �?  �>  �=  �<  �;  �:  �9  �8  �7  �6  �5  �4  �3  �2  �1  �0  �/  �.  �-  �,  �+  �*  �)  �(  �'  �&  �%  �$  �#  �"  �!  �   �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �
  �	  �  �  �  �  �  �  �  �  �   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ¾  ¼  º  ¸  ¶  ´  ²  °  ®  ¬  ª  ¨  ¦  ¤  ¢                                     �|  �x  �t  �p  �l  �h  �d  �`  �\  �X  �T  �P  �L  �H  �D  �@  �<  �8  �4  �0  �,  �(  �$  �   �  �  �  �  �  �  �  �   ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �p  �`  �P  �@  �0  �   �  �   ��  ��  ��  ��  �@  �   ��      ?�  @   @@  @�  @�  @�  @�  A   A  A   A0  A@  AP  A`  Ap  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  B   B  B  B  B  B  B  B  B   B$  B(  B,  B0  B4  B8  B<  B@  BD  BH  BL  BP  BT  BX  B\  B`  Bd  Bh  Bl  Bp  Bt  Bx  B|  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  C   C  C  C  C  C  C  C  C  C	  C
  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C   C!  C"  C#  C$  C%  C&  C'  C(  C)  C*  C+  C,  C-  C.  C/  C0  C1  C2  C3  C4  C5  C6  C7  C8  C9  C:  C;  C<  C=  C>  C?  C@  CA  CB  CC  CD  CE  CF  CG  CH  CI  CJ  CK  CL  CM  CN  CO  CP  CQ  CR  CS  CT  CU  CV  CW  CX  CY  CZ  C[  C\  C]  C^  C_  C`  Ca  Cb  Cc  Cd  Ce  Cf  Cg  Ch  Ci  Cj  Ck  Cl  Cm  Cn  Co  Cp  Cq  Cr  Cs  Ct  Cu  Cv  Cw  Cx  Cy  Cz  C{  C|  C}  C~  C  C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C�� C�  C��        	    DCAT|Waveforms|Cylinder Area   m2   UWaveform array representing the cylinder area at each point in the sample resolution. �     	   @ ����      �<-d<-$<-3e<-d<-�L<-��<.j�<.�7</z�<0�<0�n<1�O<2� <3p�<4t<5��<6�<7�<99I<:��<<=<=�.<?�<@�<Bw�<D=�<F�<G��<I�,<K�<<N�<P6�<Rk�<T��<W�<YbQ<[Ф<^L�<`��<cl<f�<h�<ky7<n@<q@<s�i<v�9<y�M<|�V<��<�l�<���<���<��<���<�P�<���<��l<�8<��<��<�9�<��<<���<�Q9<��<��t<�x�<�3�<��:<���<�i3<�'<��V<���<�b9<� �<��x<���<�X�<��<�Ͼ<���<�B.<��K<���<�b�<�z<��W<�r<�j<��_<�l�<�|<˱b<�O^<��L<Ђ<��<ӧ�<�5r<ֿ�<�F
<�ȿ<�G�<�<�9z<߬T<�<�u<��<�M]<檷<��<�W�<꧎<��<�8�<�z�<�O<��D<�"]<�P�<�y�<��<��G<�ׂ<��<���<��<��<�e<�	�<� j<��= n�= �K=S=�V=,�=��=�P=`=�7=�={�=��=+�=�=�=�=l=��=��=A=��=��=��=8�=o�=��=��=	f=	3f=	]�=	��=	��=	͎=	�=
+=
&=
>|=
TJ=
g�=
x2=
�L=
��=
��=
�6=
�=
�V=
�=
�6=
��=
��=
�K=
x2=
g�=
TJ=
>|=
&=
+=	�=	͎=	��=	��=	]�=	3f=	f=��=��=o�=8�=��=��=��=A=��=��=l=�=�=�=+�=��={�=�=�7=`=�P=��=,�=�V=S= �J= n�<��<� j<�	�<�e<��<��<���<��<�ׁ<��I<��<�y�<�P�<�"Y<��E<�O<�z�<�8�<��<꧎<�W�<��<檵<�M^<��<�u<�<߬T<�9|<�<�G�<�ȿ<�F<ֿ�<�5r<ӧ�<��<Ђ<��N<�O^<˱b<�|<�l�<��_<�j<�r<��U<�z<�b�<���<��K<�B,<���<�Ͼ<��<�X�<���<��z<� �<�b7<���<��T<�'<�i3<���<��:<�3~<�x�<��v<��<�Q9<���<��><�9�<��<��<�8<��l<���<�P�<���<��<���<���<�l�<��<|�Y<y�M<v�6<s�i<q=<n@<ky7<h�<f�<ck�<`��<^L�<[Ф<YbN<W�<T��<Rk�<P6�<N�<K�<<I�,<G��<F�<D=�<Bw�<@�<?�<=�.<<:<:��<99I<7�<6�<5��<4t<3p�<2�<1�O<0�n<0�</z�<.�7<.j�<-��<-�L<-d<-3e<-$<-d<-$<-3e<-d<-�L<-��<.j�<.�7</z�<0�<0�n<1�O<2� <3p�<4t<5��<6�<7�<99I<:��<<=<=�.<?�<@�<Bw�<D=�<F�<G��<I�,<K�<<N�<P6�<Rk�<T��<W�<YbQ<[Ф<^L�<`��<cl<f�<h�<ky7<n@<q@<s�i<v�9<y�M<|�V<��<�l�<���<���<��<���<�P�<���<��l<�8<��<��<�9�<��<<���<�Q9<��<��t<�x�<�3�<��:<���<�i3<�'<��V<���<�b9<� �<��x<���<�X�<��<�Ͼ<���<�B.<��K<���<�b�<�z<��W<�r<�j<��_<�l�<�|<˱b<�O^<��L<Ђ<��<ӧ�<�5r<ֿ�<�F
<�ȿ<�G�<�<�9z<߬T<�<�u<��<�M]<檷<��<�W�<꧎<��<�8�<�z�<�O<��D<�"]<�P�<�y�<��<��G<�ׂ<��<���<��<��<�e<�	�<� j<��= n�= �K=S=�V=,�=��=�P=`=�7=�={�=��=+�=�=�=�=l=��=��=A=��=��=��=8�=o�=��=��=	f=	3f=	]�=	��=	��=	͎=	�=
+=
&=
>|=
TJ=
g�=
x2=
�L=
��=
��=
�6=
�=
�V=
�=
�6=
��=
��=
�K=
x2=
g�=
TJ=
>|=
&=
+=	�=	͎=	��=	��=	]�=	3f=	f=��=��=o�=8�=��=��=��=A=��=��=l=�=�=�=+�=��={�=�=�7=`=�P=��=,�=�V=S= �J= n�<��<� j<�	�<�e<��<��<���<��<�ׁ<��I<��<�y�<�P�<�"Y<��E<�O<�z�<�8�<��<꧎<�W�<��<檵<�M^<��<�u<�<߬T<�9|<�<�G�<�ȿ<�F<ֿ�<�5r<ӧ�<��<Ђ<��N<�O^<˱b<�|<�l�<��_<�j<�r<��U<�z<�b�<���<��K<�B,<���<�Ͼ<��<�X�<���<��z<� �<�b7<���<��T<�'<�i3<���<��:<�3~<�x�<��v<��<�Q9<���<��><�9�<��<��<�8<��l<���<�P�<���<��<���<���<�l�<��<|�Y<y�M<v�6<s�i<q=<n@<ky7<h�<f�<ck�<`��<^L�<[Ф<YbN<W�<T��<Rk�<P6�<N�<K�<<I�,<G��<F�<D=�<Bw�<@�<?�<=�.<<:<:��<99I<7�<6�<5��<4t<3p�<2�<1�O<0�n<0�</z�<.�7<.j�<-��<-�L<-d<-3e<-$       	    DCAT|Waveforms|Exhaust Cam       eWaveform array representing the exhaust cam at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    !DCAT|Waveforms|Fuel Rail Pressure   MPa   lWaveform array representing the fuel rail pressure at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|HRR   J/CAD   kWaveform array representing the heat release rate at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Injector Command       jWaveform array representing the injector command at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    "DCAT|Waveforms|Instantaneous Speed   RPM   mWaveform array representing the instantaneous speed at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Intake Cam       dWaveform array representing the intake cam at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|MFB   Fraction   nWaveform array representing the mass fraction burned at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    )DCAT|Waveforms|Manifold Absolute Pressure   kPa abs   tWaveform array representing the manifold absolute pressure at each point in the sample resolution for each cylinder. �     	   @ ��������                     
     DCAT|Waveforms|Motoring Pressure   kPa abs   kWaveform array representing the Motoring pressure at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|PWM       �Waveform array representing the pulse width modulation at each point in the sample resolution for each cylinder. The data is stored in a bitfield representing each pulse width modulation channel. �     	   @ ��������                     
    DCAT|Waveforms|PWM Names       ZName or description associated with each pulse width modulation channel and each cylinder. �     0����                  "DCAT|Waveforms|PreChamber Pressure   kPa abs   nWaveform array representing the pre chamber pressure at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Pressure   kPa abs   kWaveform array representing the cylinder pressure at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Spark Command       gWaveform array representing the spark command at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Synchronous Pump       jWaveform array representing the synchronous pump at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|TDC Probe       oWaveform array representing the top dead center probe at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Temp   K   rWaveform array representing the cylinder gas temperature at each point in the sample resolution for each cylinder. �     	   @ ��������                     
    DCAT|Waveforms|Volume   liter   YWaveform array representing the calculated volume at each point in the sample resolution. �     	   @ ����      �<�<�j<��<��W<�D&<��R<��= �=��=EK=	�=d=t2=E?=v="='�g=.@^=4�%=;��=CM�=K�=S�=[�(=dHz=m`�=v��=�GR=�P�=�� =��=�^V=�)=���=�Ə=�ݶ=�j=�v=���=Ɩ�=�W�=�8�=�8d=�U�=鐌=��D=�YI=��>ź>��>��>�A>�s>�>��>Ǧ>#�>( >,X�>0��>4߹>9-`>=�>Aځ>F9>J�*>O>Sn�>W��>\M�>`�E>e6w>i�>n$�>r��>w�>{�1>�|>�<A>�v)>��>��>��>�Q<>���>��m>���>��>�8>�^�>��#>���>���>�ْ>��>�">��>� >�!j>�#f>� �>��>�/>���>��3>�͵>��>��>>�_>�/p>��O>ſ�>�->�9>��>̛ >�CF>��d>сm>�P>ԧ>�0y>׳�>�0u>ڦ�>��>݀�>��>�@S>�i>���>�.�>�q@>��>��>��>�8S>�Yp>�s�>퇛>>��>�>�>��>�qK>�V>�4.>��>��<>��4>�ix>�&>���>��%>�3�>�Պ>�p�>�?>��>�V>���>��>��'>���? -r? ],? ��? ��? ؈? �?H?69?N�?d8?vJ?�?��?��?��?�X?��?��?��?�?vI?d8?N�?69?H? �? ؈? ��? ��? ],? -r>���>��'>��>���>�V>��>�?>�p�>�Պ>�3�>��%>���>�&>�iz>��4>��:>��>�4.>�V>�qK>��>�>�>� >>퇝>�s�>�Yp>�8Q>��>��>��>�q@>�.�>���>�i>�@P>��>݀�>��>ڦ�>�0u>׳�>�0u>ԧ>�P>сk>��b>�CF>̛ >��>�9>�+>ſ�>��O>�/p>�_>��>>��>�͵>��1>���>�->��>� �>�#f>�!j>�>��>�">��>�ْ>���>���>��#>�^�>�7�>��>���>��m>���>�Q:>��>��>��>�v)>�<A>�~>{�5>w�>r��>n$�>i�>e6w>`�E>\M�>W��>Sn�>O�>J�*>F9>A�}>=�">9-`>4߹>0��>,X�>( >#�>Ǣ>��>�>�s>�=>��>��>ž=��=�YA=��D=鐃=�U�=�8d=�8�=�W�=Ɩ�=���=�v=�j=�ݮ=�Ə=���=�)=�^V=��=�� =�P�=�GR=v��=m`�=dHz=[�(=S�=K�=CM�=;��=4�%=.@^='�g="=v=E?=t!=d=	�=EK=��= �<��<��0<�D&<��W<��<�j<�<�j<��<��W<�D&<��R<��= �=��=EK=	�=d=t2=E?=v="='�g=.@^=4�%=;��=CM�=K�=S�=[�(=dHz=m`�=v��=�GR=�P�=�� =��=�^V=�)=���=�Ə=�ݶ=�j=�v=���=Ɩ�=�W�=�8�=�8d=�U�=鐌=��D=�YI=��>ź>��>��>�A>�s>�>��>Ǧ>#�>( >,X�>0��>4߹>9-`>=�>Aځ>F9>J�*>O>Sn�>W��>\M�>`�E>e6w>i�>n$�>r��>w�>{�1>�|>�<A>�v)>��>��>��>�Q<>���>��m>���>��>�8>�^�>��#>���>���>�ْ>��>�">��>� >�!j>�#f>� �>��>�/>���>��3>�͵>��>��>>�_>�/p>��O>ſ�>�->�9>��>̛ >�CF>��d>сm>�P>ԧ>�0y>׳�>�0u>ڦ�>��>݀�>��>�@S>�i>���>�.�>�q@>��>��>��>�8S>�Yp>�s�>퇛>>��>�>�>��>�qK>�V>�4.>��>��<>��4>�ix>�&>���>��%>�3�>�Պ>�p�>�?>��>�V>���>��>��'>���? -r? ],? ��? ��? ؈? �?H?69?N�?d8?vJ?�?��?��?��?�X?��?��?��?�?vI?d8?N�?69?H? �? ؈? ��? ��? ],? -r>���>��'>��>���>�V>��>�?>�p�>�Պ>�3�>��%>���>�&>�iz>��4>��:>��>�4.>�V>�qK>��>�>�>� >>퇝>�s�>�Yp>�8Q>��>��>��>�q@>�.�>���>�i>�@P>��>݀�>��>ڦ�>�0u>׳�>�0u>ԧ>�P>сk>��b>�CF>̛ >��>�9>�+>ſ�>��O>�/p>�_>��>>��>�͵>��1>���>�->��>� �>�#f>�!j>�>��>�">��>�ْ>���>���>��#>�^�>�7�>��>���>��m>���>�Q:>��>��>��>�v)>�<A>�~>{�5>w�>r��>n$�>i�>e6w>`�E>\M�>W��>Sn�>O�>J�*>F9>A�}>=�">9-`>4߹>0��>,X�>( >#�>Ǣ>��>�>�s>�=>��>��>ž=��=�YA=��D=鐃=�U�=�8d=�8�=�W�=Ɩ�=���=�v=�j=�ݮ=�Ə=���=�)=�^V=��=�� =�P�=�GR=v��=m`�=dHz=[�(=S�=K�=CM�=;��=4�%=.@^='�g="=v=E?=t!=d=	�=EK=��= �<��<��0<�D&<��W<��<�j       	    DCAT|Waveforms|dVolume   liter   UWaveform array representing the volume change at each point in the sample resolution. �     	   @ ����      �8G� 8�� 9G�@9��`9ǟ`9�T�:s�:..�:F�`:_X�:w� :�	 :��:�0:��:�� :ä :�K�:��@:�J :�`:�� ;�;	m;��;+p;n ;�P;#��;(�p;-�`;2��;7W;<`;@��;E�;I��;M�`;R�;V#;Z#;^	0;a��;e��;i�;l��;o�;s"�;vC�;yF@;|*�;~��;�� ;��;�I0;�o�;��@;��;���;�r�;�K�;�P;��;�~�;��;���;�&P;���;���;�F�;���;��p;��;��`;� @;���;�� ;��;���;�X`;��;���;�S�;��`;�f ;���;�H ;�� ;���;�D ;�� ;�� ;���;���;� ;��;��;��;��;��;}� ;{P�;x�@;v� ;t�;qy ;n�@;l=�;i��;f�@;d@;a7�;^\@;[u�;X��;U��;R� ;O��;L{ ;Ie ;FJ@;C'�;?� ;<��;9�@;6j ;3/@;/�@;,��;)g�;& ;"��;��;5�;��;�@;:�;� ;��;1�;��;@:�I :�� :�݀:�'�:�q�:ڼ :� :�S :ƞ :��:�=�:�� :�� :�2�:���:�ڀ:�2 :���:��:z� :m> :`  :R� :E� :8J :+ :� :� :� 9� 9�P 9�� 9�� 9�h 9R( 9� 8�P 8R@     �R@ ��P �� �R0 ��h ��� ��� ��P �� �� �� �� �+ �8J �E� �R� �`  �m> �z� ��怺�����2 ��ڀ������2���� ��� ��<���퀺Ơ ��S �� �ڼ ��q���'���݀��� ��H �@����1���@�〻: �����@�5�����"���& �)h@�,���/� �3.��6i��9���<���@  �C' �FI@�If �L{��O�@�R���U���X���[v �^[��a7 �d��f���i���l<��n�@�qz �t��v� �x�@�{P �}� �����	 ��`�����໅ ��� ����������� ��D�����������H ��� ��f`���`��S����������X`���`���л�栻��p�� @��� ���p���p���໎Fໍ�����@��&P���л�л�~@���л����L��r@���P����������oໃH������͠�~��|*��yE��vC@�s#��o倻l��i �e��a��^	0�Z#�V"��R �M��I�0�E��@��<`�7W��2���-�`�(�p�#���P�n��+p��@�	m������`��I���@��K�ä ��� ��к�@������w� �_X��F�`�..�v ��T��Ǜ ���`�G�@��8G� 8�� 9G�@9��`9ǟ`9�T�:s�:..�:F�`:_X�:w� :�	 :��:�0:��:�� :ä :�K�:��@:�J :�`:�� ;�;	m;��;+p;n ;�P;#��;(�p;-�`;2��;7W;<`;@��;E�;I��;M�`;R�;V#;Z#;^	0;a��;e��;i�;l��;o�;s"�;vC�;yF@;|*�;~��;�� ;��;�I0;�o�;��@;��;���;�r�;�K�;�P;��;�~�;��;���;�&P;���;���;�F�;���;��p;��;��`;� @;���;�� ;��;���;�X`;��;���;�S�;��`;�f ;���;�H ;�� ;���;�D ;�� ;�� ;���;���;� ;��;��;��;��;��;}� ;{P�;x�@;v� ;t�;qy ;n�@;l=�;i��;f�@;d@;a7�;^\@;[u�;X��;U��;R� ;O��;L{ ;Ie ;FJ@;C'�;?� ;<��;9�@;6j ;3/@;/�@;,��;)g�;& ;"��;��;5�;��;�@;:�;� ;��;1�;��;@:�I :�� :�݀:�'�:�q�:ڼ :� :�S :ƞ :��:�=�:�� :�� :�2�:���:�ڀ:�2 :���:��:z� :m> :`  :R� :E� :8J :+ :� :� :� 9� 9�P 9�� 9�� 9�h 9R( 9� 8�P 8R@     �R@ ��P �� �R0 ��h ��� ��� ��P �� �� �� �� �+ �8J �E� �R� �`  �m> �z� ��怺�����2 ��ڀ������2���� ��� ��<���퀺Ơ ��S �� �ڼ ��q���'���݀��� ��H �@����1���@�〻: �����@�5�����"���& �)h@�,���/� �3.��6i��9���<���@  �C' �FI@�If �L{��O�@�R���U���X���[v �^[��a7 �d��f���i���l<��n�@�qz �t��v� �x�@�{P �}� �����	 ��`�����໅ ��� ����������� ��D�����������H ��� ��f`���`��S����������X`���`���л�栻��p�� @��� ���p���p���໎Fໍ�����@��&P���л�л�~@���л����L��r@���P����������oໃH������͠�~��|*��yE��vC@�s#��o倻l��i �e��a��^	0�Z#�V"��R �M��I�0�E��@��<`�7W��2���-�`�(�p�#���P�n��+p��@�	m������`��I���@��K�ä ��� ��к�@������w� �_X��F�`�..�v ��T��Ǜ ���`�G�@��       	    D|Fuel|ClosedLoopDieselFuelOn   |   .Indicated is closed loop fuel contro is active �     !               ECS|ADCombo|ADComboPresent   |   0Indicates AD Combo module's presence is detected �     !              ECS|Boost|Boost1ControlKp       Boost PID Kp �     	                  ECS|Boost|Boost1ControlTd   min   Boost PID Td �     	                  ECS|Boost|Boost1ControlTi   min   Boost PID Ti �     	                  ECS|Boost|Boost1DC   %   Final Boost Duty Cycle �     	                   ECS|Boost|Boost1Enable   |     �     !              ECS|Boost|Boost1Freq         �     	                  ECS|Boost|Boost1PIDEnable   |   Enable Boost PID �     !              ECS|Boost|Boost1Setpoint   bar   Boost PID Setpoint �     	    ?�             ECS|Boost|Boost1Table   mm3/cyc|rpm|bar   Boost Pressure Setpoint Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  A   A   AP  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ� Ej` Ez  E�� E�� E�p E�@       ?�  ?�  ?�G�?��\?��?���?�33?���?�  ?�ff?���?�33?���?��H?�  ?�  ?�  ?�%?�33?�?��?��?�Q�?�{?�z�?��H?�%?�
=?�(�?���?�9X?�9X?�  ?��?��?�ff?�=q?�
=?�p�?��\?���?�\)?��?��H?��R?�M�?�Q�?�Q�?�G�?��
?�?�ff?���?���?���?�Q�?��R?�E�?���?���?���?�r�?͑h?̋D?��/?�l�?�ff?���?�
=?���?��^?�{?�z�?�/?�M�?�Q�?�C�?Η�?ҏ\?У�?���?���?���?�?�(�?���?�S�?�l�?�p�?öF?���?�v�?�n�?�?�b?��?���?�{?��?��?�G�?�
=?��H?�\)?�z�?�=q?�\)?�z�?ٙ�?�p�?�p�?�33?�%?�\)?�
=?�G�?�=q?�(�?öF?�=q?��m?�hs?�ff?ۅ?�  ?�S�?��?��
?��?�?�p�?�ff?�z�?�?̋D?��
?�?ش9?�p�?�\?�ff?�X?�ff?�z�?�  ?�l�?�\)?�
=?���?�
=?�(�?�33?��
?�
=?陚?�|�?�\?�?�Ĝ?�z�?���?�ff?�  ?�{?׮?��T?陚?�G�?��?�z�?��?�{@   @   ?���?�z�?��
?�  ?���?�{?陚?�33?�@   @G�@33@@\)@ff@ff@�?�z�?��?Ǯ?�(�?���@   @�
@ff@\)@"�@1@�@��@��@p�@
�H?�z�?��?�z�?��@ff@
J@�@(�@{@z�@@ff@
=@��@p�@
�H?�z�?��?�  ?�(�@Q�@p�@��@=q@z�@�@@ff@
=@��@p�@
�H?�z�?��?�  @�@	��@p�@��@=q@z�@�@@ff@
=@��@p�@
�H?�z�          ECS|Boost|Boost2ControlKp       Boost PID Kp �     	                  ECS|Boost|Boost2ControlTd   min   Boost PID Td �     	                  ECS|Boost|Boost2ControlTi   min   Boost PID Ti �     	                  ECS|Boost|Boost2DC   %   Final Boost Duty Cycle �     	                   ECS|Boost|Boost2Enable   |     �     !              ECS|Boost|Boost2Freq         �     	                  ECS|Boost|Boost2PIDEnable   |   Enable Boost PID �     !              ECS|Boost|Boost2Setpoint   bar   Boost PID Setpoint �     	    ?�             ECS|Boost|Boost2Table   mm3/cyc|rpm|bar   Boost Pressure Setpoint Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  A   A   AP  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ� Ej` Ez  E�� E�� E�p E�@       ?�  ?�  ?�G�?��\?��?���?�33?���?�  ?�ff?���?�33?���?��H?�  ?�  ?�  ?�%?�33?�?��?��?�Q�?�{?�z�?��H?�%?�
=?�(�?���?�9X?�9X?�  ?��?��?�ff?�=q?�
=?�p�?��\?���?�\)?��?��H?��R?�M�?�Q�?�Q�?�G�?��
?�?�ff?���?���?���?�Q�?��R?�E�?���?���?���?�r�?͑h?̋D?��/?�l�?�ff?���?�
=?���?��^?�{?�z�?�/?�M�?�Q�?�C�?Η�?ҏ\?У�?���?���?���?�?�(�?���?�S�?�l�?�p�?öF?���?�v�?�n�?�?�b?��?���?�{?��?��?�G�?�
=?��H?�\)?�z�?�=q?�\)?�z�?ٙ�?�p�?�p�?�33?�%?�\)?�
=?�G�?�=q?�(�?öF?�=q?��m?�hs?�ff?ۅ?�  ?�S�?��?��
?��?�?�p�?�ff?�z�?�?̋D?��
?�?ش9?�p�?�\?�ff?�X?�ff?�z�?�  ?�l�?�\)?�
=?���?�
=?�(�?�33?��
?�
=?陚?�|�?�\?�?�Ĝ?�z�?���?�ff?�  ?�{?׮?��T?陚?�G�?��?�z�?��?�{@   @   ?���?�z�?��
?�  ?���?�{?陚?�33?�@   @G�@33@@\)@ff@ff@�?�z�?��?Ǯ?�(�?���@   @�
@ff@\)@"�@1@�@��@��@p�@
�H?�z�?��?�z�?��@ff@
J@�@(�@{@z�@@ff@
=@��@p�@
�H?�z�?��?�  ?�(�@Q�@p�@��@=q@z�@�@@ff@
=@��@p�@
�H?�z�?��?�  @�@	��@p�@��@=q@z�@�@@ff@
=@��@p�@
�H?�z�          ECS|Boost|DesBoost1DC   %   .Desired Boost Duty Cycle before Manual Setting �     	                   ECS|Boost|DesBoost1Setpoint   bar   ,Desired Boost Setpoint before Manual Setting �     	    ?�             ECS|Boost|DesBoost2DC   %   .Desired Boost Duty Cycle before Manual Setting �     	                   ECS|Boost|DesBoost2Setpoint   bar   ,Desired Boost Setpoint before Manual Setting �     	    ?�             ECS|Boost|DesWGDC   %   .Desired Boost Duty Cycle before Manual Setting �     	                   ECS|Boost|DesWGSetpoint   bar   ,Desired Boost Setpoint before Manual Setting �     	    ?�             ECS|Boost|ManualBoost1DC   %   Manual Boost Duty Cycle Setting �     	                  ECS|Boost|ManualBoost1DCEnable   Manual|Automatic   -Override boost duty cycle with manual setting �     !              ECS|Boost|ManualBoost1Setpoint   bar   Manual Boost Setting �     	                  $ECS|Boost|ManualBoost1SetpointEnable   Manual|Automatic   +Override boost setpoint with manual setting �     !              ECS|Boost|ManualBoost2DC   %   Manual Boost Duty Cycle Setting �     	                  ECS|Boost|ManualBoost2DCEnable   Manual|Automatic   -Override boost duty cycle with manual setting �     !              ECS|Boost|ManualBoost2Setpoint   bar   Manual Boost Setting �     	                  $ECS|Boost|ManualBoost2SetpointEnable   Manual|Automatic   +Override boost setpoint with manual setting �     !              ECS|Boost|ManualWGDC   %   Manual Boost Duty Cycle Setting �     	                  ECS|Boost|ManualWGDCEnable   Manual|Automatic   -Override boost duty cycle with manual setting �     !              ECS|Boost|ManualWGSetpoint   bar   Manual Boost Setting �     	                   ECS|Boost|ManualWGSetpointEnable   Manual|Automatic   +Override boost setpoint with manual setting �     !              ECS|Boost|MaxBoost1DC   %   Max Boost Duty Cycle �     	                  ECS|Boost|MaxBoost2DC   %   Max Boost Duty Cycle �     	                  ECS|Boost|MaxWGDC   %   Max Boost Duty Cycle �     	                  ECS|Boost|MinBoost1DC   %   Min Boost Duty Cycle �     	                  ECS|Boost|MinBoost2DC   %   Min Boost Duty Cycle �     	                  ECS|Boost|MinWGDC   %   Min Boost Duty Cycle �     	                  ECS|Boost|WGControlKp       Boost PID Kp �     	                  ECS|Boost|WGControlTd   min   Boost PID Td �     	                  ECS|Boost|WGControlTi   min   Boost PID Ti �     	                  ECS|Boost|WGDC   %   Final Boost Duty Cycle �     	                   ECS|Boost|WGPIDEnable   |   Enable Boost PID �     !              ECS|Boost|WGSetpoint   bar   Boost PID Setpoint �     	    ?�             ECS|Boost|WGTable   mm3/cyc|rpm|bar   Boost Pressure Setpoint Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  A   A   AP  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ� Ej` Ez  E�� E�� E�p E�@       ?�  ?�  ?�G�?��\?��?���?�33?���?�  ?�ff?���?�33?���?��H?�  ?�  ?�  ?�%?�33?�?��?��?�Q�?�{?�z�?��H?�%?�
=?�(�?���?�9X?�9X?�  ?��?��?�ff?�=q?�
=?�p�?��\?���?�\)?��?��H?��R?�M�?�Q�?�Q�?�G�?��
?�?�ff?���?���?���?�Q�?��R?�E�?���?���?���?�r�?͑h?̋D?��/?�l�?�ff?���?�
=?���?��^?�{?�z�?�/?�M�?�Q�?�C�?Η�?ҏ\?У�?���?���?���?�?�(�?���?�S�?�l�?�p�?öF?���?�v�?�n�?�?�b?��?���?�{?��?��?�G�?�
=?��H?�\)?�z�?�=q?�\)?�z�?ٙ�?�p�?�p�?�33?�%?�\)?�
=?�G�?�=q?�(�?öF?�=q?��m?�hs?�ff?ۅ?�  ?�S�?��?��
?��?�?�p�?�ff?�z�?�?̋D?��
?�?ش9?�p�?�\?�ff?�X?�ff?�z�?�  ?�l�?�\)?�
=?���?�
=?�(�?�33?��
?�
=?陚?�|�?�\?�?�Ĝ?�z�?���?�ff?�  ?�{?׮?��T?陚?�G�?��?�z�?��?�{@   @   ?���?�z�?��
?�  ?���?�{?陚?�33?�@   @G�@33@@\)@ff@ff@�?�z�?��?Ǯ?�(�?���@   @�
@ff@\)@"�@1@�@��@��@p�@
�H?�z�?��?�z�?��@ff@
J@�@(�@{@z�@@ff@
=@��@p�@
�H?�z�?��?�  ?�(�@Q�@p�@��@=q@z�@�@@ff@
=@��@p�@
�H?�z�?��?�  @�@	��@p�@��@=q@z�@�@@ff@
=@��@p�@
�H?�z�          ECS|CriticalFault|FPGA_1_Error   Failed|Success   1Indicates FPGA did not load.  Recompile required. �     !               ECS|CriticalFault|FPGA_2_Error   Failed|Success   1Indicates FPGA did not load.  Recompile required. �     !               ECS|DI1|DI1_BackBoostTime   msec   xTime period during which injector solenoid energy is directed back to the module boost power supply (after end of pulse) �     	    >��          ECS|DI1|DI1_BatteryVoltage       DI Driver battery voltage level �     	                   ECS|DI1|DI1_Chan1Enable   |   "Enables channel regardless of mode �     !             ECS|DI1|DI1_Chan2Enable   |   "Enables channel regardless of mode �     !             ECS|DI1|DI1_ClearFaults   ON|OFF   )Clears any critical faults with DI Driver �     !              ECS|DI1|DI1_ExternalHighVoltage       cHigh voltage level supplied externally to terminal 7 of DI Driver to override internal boost supply �     	                   ECS|DI1|DI1_FI1OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI1|DI1_FI2OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI1|DI1_FI3OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI1|DI1_HVTarget   V   9DI Driver high voltage setpoint for internal boost supply �     	    B�            "ECS|DI1|DI1_HighVoltageDriverFault   FAULT|NO FAULT   !High voltage driver circuit fault �     !               !ECS|DI1|DI1_HighVoltageLimitFault   FAULT|NO FAULT   .Internal boost power supply over-voltage fault �     !               ECS|DI1|DI1_InjectionEnable   ON|OFF   Enables all channels of module �     !             ECS|DI1|DI1_InternalHighVoltage       (Internal boost supply high voltage level �     	                   !ECS|DI1|DI1_LowVoltageDriverFault   FAULT|NO FAULT    Low voltage driver circuit fault �     !               ECS|DI1|DI1_ModuleEnable   ON|OFF   "Enables DI Driver module operation �     !              ECS|DI1|DI1_ModulePresent   ON|OFF   9Indicates DI Driver module present and externally powered �     !               ECS|DI1|DI1_ModuleRev       0Indicates DI Driver module Hardware/Firmware Rev �     0����                  ECS|DI1|DI1_ModuleTempFault   FAULT|NO FAULT   #Module over-temperature fault (80C) �     !               ECS|DI1|DI1_ModuleTemperature       Internal module temperature �     	                   ECS|DI1|DI1_OLIntegrator       3Indicates level of internal boost power supply load �                        ECS|DI1|DI1_OneShot   FIRE NOW|OFF   .Generates one-shot command to selected channel �     !              ECS|DI1|DI1_OneShotSelect   Disabled|Chan 1|Chan 2|Chan 3   $Selects channel for one-shot command �                      ECS|DI1|DI1_OneShotTime   msec   Duration of one-shot command �     	    ?�            ECS|DI1|DI1_OpenCircuitOverride   ON|OFF   4Determines whether open-circuit faults are indicated �     !              ECS|DI1|DI1_PSChargeFault   FAULT|NO FAULT   *Internal boost power supply charging fault �     !               ECS|DI1|DI1_PSOverloadFault   FAULT|NO FAULT   *Internal boost power supply overload fault �     !               !ECS|DI1|DI1_Phase1FirstPeakEnable   ON|OFF   8Causes phase 2 to begin after current reaches first peak �     !             ECS|DI1|DI1_PiezoEnable   ON|OFF   Enables piezo operating mode �     !              ECS|DI1|DI1_PiezoInvert   ON|OFF   %Enables inverted piezo operating mode �     !              ECS|DI1|DI1_PowerSupplyEnable   ON|OFF   #Enables internal boost power supply �     !             ECS|DI1|DI1_ShortCircuitFault   FAULT|NO FAULT   Injector short-circuit fault �     !               ECS|DI2|DI2_BackBoostTime   msec   xTime period during which injector solenoid energy is directed back to the module boost power supply (after end of pulse) �     	    >��          ECS|DI2|DI2_BatteryVoltage       DI Driver battery voltage level �     	                   ECS|DI2|DI2_Chan1Enable   |   "Enables channel regardless of mode �     !              ECS|DI2|DI2_Chan2Enable   |   "Enables channel regardless of mode �     !              ECS|DI2|DI2_ClearFaults   ON|OFF   )Clears any critical faults with DI Driver �     !              ECS|DI2|DI2_ExternalHighVoltage       cHigh voltage level supplied externally to terminal 7 of DI Driver to override internal boost supply �     	                   ECS|DI2|DI2_FI1OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI2|DI2_FI2OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI2|DI2_FI3OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI2|DI2_HVTarget   V   9DI Driver high voltage setpoint for internal boost supply �     	    B�            "ECS|DI2|DI2_HighVoltageDriverFault   FAULT|NO FAULT   !High voltage driver circuit fault �     !               !ECS|DI2|DI2_HighVoltageLimitFault   FAULT|NO FAULT   .Internal boost power supply over-voltage fault �     !               ECS|DI2|DI2_InjectionEnable   ON|OFF   Enables all channels of module �     !              ECS|DI2|DI2_InternalHighVoltage       (Internal boost supply high voltage level �     	                   !ECS|DI2|DI2_LowVoltageDriverFault   FAULT|NO FAULT    Low voltage driver circuit fault �     !               ECS|DI2|DI2_ModuleEnable   ON|OFF   "Enables DI Driver module operation �     !              ECS|DI2|DI2_ModulePresent   ON|OFF   9Indicates DI Driver module present and externally powered �     !               ECS|DI2|DI2_ModuleRev       0Indicates DI Driver module Hardware/Firmware Rev �     0����                  ECS|DI2|DI2_ModuleTempFault   FAULT|NO FAULT   #Module over-temperature fault (80C) �     !               ECS|DI2|DI2_ModuleTemperature       Internal module temperature �     	                   ECS|DI2|DI2_OLIntegrator       3Indicates level of internal boost power supply load �                        ECS|DI2|DI2_OneShot   FIRE NOW|OFF   .Generates one-shot command to selected channel �     !              ECS|DI2|DI2_OneShotSelect   Disabled|Chan 1|Chan 2|Chan 3   $Selects channel for one-shot command �                       ECS|DI2|DI2_OneShotTime   msec   Duration of one-shot command �     	    ?�            ECS|DI2|DI2_OpenCircuitOverride   ON|OFF   4Determines whether open-circuit faults are indicated �     !              ECS|DI2|DI2_PSChargeFault   FAULT|NO FAULT   *Internal boost power supply charging fault �     !               ECS|DI2|DI2_PSOverloadFault   FAULT|NO FAULT   *Internal boost power supply overload fault �     !               !ECS|DI2|DI2_Phase1FirstPeakEnable   ON|OFF   8Causes phase 2 to begin after current reaches first peak �     !              ECS|DI2|DI2_PiezoEnable   ON|OFF   Enables piezo operating mode �     !              ECS|DI2|DI2_PiezoInvert   ON|OFF   %Enables inverted piezo operating mode �     !              ECS|DI2|DI2_PowerSupplyEnable   ON|OFF   #Enables internal boost power supply �     !              ECS|DI2|DI2_ShortCircuitFault   FAULT|NO FAULT   Injector short-circuit fault �     !               ECS|DI3|DI3_BackBoostTime   msec   xTime period during which injector solenoid energy is directed back to the module boost power supply (after end of pulse) �     	    >��          ECS|DI3|DI3_BatteryVoltage       DI Driver battery voltage level �     	                   ECS|DI3|DI3_Chan1Enable   |   "Enables channel regardless of mode �     !              ECS|DI3|DI3_Chan2Enable   |   "Enables channel regardless of mode �     !              ECS|DI3|DI3_ClearFaults   ON|OFF   )Clears any critical faults with DI Driver �     !              ECS|DI3|DI3_ExternalHighVoltage       cHigh voltage level supplied externally to terminal 7 of DI Driver to override internal boost supply �     	                   ECS|DI3|DI3_FI1OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI3|DI3_FI2OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI3|DI3_FI3OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI3|DI3_HVTarget   V   9DI Driver high voltage setpoint for internal boost supply �     	    B�            "ECS|DI3|DI3_HighVoltageDriverFault   FAULT|NO FAULT   !High voltage driver circuit fault �     !               !ECS|DI3|DI3_HighVoltageLimitFault   FAULT|NO FAULT   .Internal boost power supply over-voltage fault �     !               ECS|DI3|DI3_InjectionEnable   ON|OFF   Enables all channels of module �     !              ECS|DI3|DI3_InternalHighVoltage       (Internal boost supply high voltage level �     	                   !ECS|DI3|DI3_LowVoltageDriverFault   FAULT|NO FAULT    Low voltage driver circuit fault �     !               ECS|DI3|DI3_ModuleEnable   ON|OFF   "Enables DI Driver module operation �     !              ECS|DI3|DI3_ModulePresent   ON|OFF   9Indicates DI Driver module present and externally powered �     !               ECS|DI3|DI3_ModuleRev       0Indicates DI Driver module Hardware/Firmware Rev �     0����                  ECS|DI3|DI3_ModuleTempFault   FAULT|NO FAULT   #Module over-temperature fault (80C) �     !               ECS|DI3|DI3_ModuleTemperature       Internal module temperature �     	                   ECS|DI3|DI3_OLIntegrator       3Indicates level of internal boost power supply load �                        ECS|DI3|DI3_OneShot   FIRE NOW|OFF   .Generates one-shot command to selected channel �     !              ECS|DI3|DI3_OneShotSelect   Disabled|Chan 1|Chan 2|Chan 3   $Selects channel for one-shot command �                       ECS|DI3|DI3_OneShotTime   msec   Duration of one-shot command �     	    ?�            ECS|DI3|DI3_OpenCircuitOverride   ON|OFF   4Determines whether open-circuit faults are indicated �     !              ECS|DI3|DI3_PSChargeFault   FAULT|NO FAULT   *Internal boost power supply charging fault �     !               ECS|DI3|DI3_PSOverloadFault   FAULT|NO FAULT   *Internal boost power supply overload fault �     !               !ECS|DI3|DI3_Phase1FirstPeakEnable   ON|OFF   8Causes phase 2 to begin after current reaches first peak �     !              ECS|DI3|DI3_PiezoEnable   ON|OFF   Enables piezo operating mode �     !              ECS|DI3|DI3_PiezoInvert   ON|OFF   %Enables inverted piezo operating mode �     !              ECS|DI3|DI3_PowerSupplyEnable   ON|OFF   #Enables internal boost power supply �     !              ECS|DI3|DI3_ShortCircuitFault   FAULT|NO FAULT   Injector short-circuit fault �     !               ECS|DI4|DI4_BackBoostTime   msec   xTime period during which injector solenoid energy is directed back to the module boost power supply (after end of pulse) �     	    >��          ECS|DI4|DI4_BatteryVoltage       DI Driver battery voltage level �     	                   ECS|DI4|DI4_Chan1Enable   |   "Enables channel regardless of mode �     !              ECS|DI4|DI4_Chan2Enable   |   "Enables channel regardless of mode �     !              ECS|DI4|DI4_ClearFaults   ON|OFF   )Clears any critical faults with DI Driver �     !              ECS|DI4|DI4_ExternalHighVoltage       cHigh voltage level supplied externally to terminal 7 of DI Driver to override internal boost supply �     	                   ECS|DI4|DI4_FI1OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI4|DI4_FI2OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI4|DI4_FI3OpenCircuit   FAULT|NO FAULT   Injector open-circuit fault �     !               ECS|DI4|DI4_HVTarget   V   9DI Driver high voltage setpoint for internal boost supply �     	    B�            "ECS|DI4|DI4_HighVoltageDriverFault   FAULT|NO FAULT   !High voltage driver circuit fault �     !               !ECS|DI4|DI4_HighVoltageLimitFault   FAULT|NO FAULT   .Internal boost power supply over-voltage fault �     !               ECS|DI4|DI4_InjectionEnable   ON|OFF   Enables all channels of module �     !              ECS|DI4|DI4_InternalHighVoltage       (Internal boost supply high voltage level �     	                   !ECS|DI4|DI4_LowVoltageDriverFault   FAULT|NO FAULT    Low voltage driver circuit fault �     !               ECS|DI4|DI4_ModuleEnable   ON|OFF   "Enables DI Driver module operation �     !              ECS|DI4|DI4_ModulePresent   ON|OFF   9Indicates DI Driver module present and externally powered �     !               ECS|DI4|DI4_ModuleRev       0Indicates DI Driver module Hardware/Firmware Rev �     0����                  ECS|DI4|DI4_ModuleTempFault   FAULT|NO FAULT   #Module over-temperature fault (80C) �     !               ECS|DI4|DI4_ModuleTemperature       Internal module temperature �     	                   ECS|DI4|DI4_OLIntegrator       3Indicates level of internal boost power supply load �                        ECS|DI4|DI4_OneShot   FIRE NOW|OFF   .Generates one-shot command to selected channel �     !              ECS|DI4|DI4_OneShotSelect   Disabled|Chan 1|Chan 2|Chan 3   $Selects channel for one-shot command �                       ECS|DI4|DI4_OneShotTime   msec   Duration of one-shot command �     	    ?�            ECS|DI4|DI4_OpenCircuitOverride   ON|OFF   4Determines whether open-circuit faults are indicated �     !              ECS|DI4|DI4_PSChargeFault   FAULT|NO FAULT   *Internal boost power supply charging fault �     !               ECS|DI4|DI4_PSOverloadFault   FAULT|NO FAULT   *Internal boost power supply overload fault �     !               !ECS|DI4|DI4_Phase1FirstPeakEnable   ON|OFF   8Causes phase 2 to begin after current reaches first peak �     !              ECS|DI4|DI4_PiezoEnable   ON|OFF   Enables piezo operating mode �     !              ECS|DI4|DI4_PiezoInvert   ON|OFF   %Enables inverted piezo operating mode �     !              ECS|DI4|DI4_PowerSupplyEnable   ON|OFF   #Enables internal boost power supply �     !              ECS|DI4|DI4_ShortCircuitFault   FAULT|NO FAULT   Injector short-circuit fault �     !               ECS|DI|DIFuelDurationArray   msec   DI Fuel Duration Array �     	   @ ����               ?�                 	    ECS|DI|DIFuelTimingArray   DBTDC   DI Fuel Timing Array �     	   @ ����       Bp  Bp      �   �          	    ECS|DI|DI_Window_End   DBTDC   Spark Operating Window Start �     	    �p            ECS|DI|DI_Window_Start   DBTDC   Spark Operating Window Start �     	    Bp            ECS|DI|IPhaseCurrentLower       iPhase Current Lower Limit �     	   @ ����       A�  A`                                 	   ECS|DI|IPhaseCurrentUpper       iPhase Current Upper Limit �     	   @ ����       A�  Ap                                 	   ECS|DI|IPhaseDrive       <Selects low voltage or high voltage for the associated phase �                    ECS|DI|IPhaseDuration       iPhase Duration �     	   @ ����       =���                                   	   ECS|DiffIO1|DiffIO1_Init   ON|OFF   .Initialize DiffIO Module for Direction Control �     !              !ECS|DiffIO1|DiffIO1_ModulePresent   ON|OFF   :Indicates PFI Driver module present and externally powered �     !              "ECS|DiffIO1|DiffIO1_ModulePresent2   ON|OFF   :Indicates PFI Driver module present and externally powered �     !               ECS|EGR|HPEGRFreq         �     	                  ECS|EGR|LPEGREnable   |     �     !              ECS|EGR|LPEGRFreq         �     	                  ECS|EGR|ThrottleFreq         �     	                  "ECS|EPT|AutoClearFlagWhileCranking   |   3Auto-clears EPT errors during EngineStatus=CRANKING �     !              ECS|EPT|Cam1_DigChanAsn_Mem       +Assigns digital signal source to cam signal �         
           ECS|EPT|Cam2_DigChanAsn_Mem       +Assigns digital signal source to cam signal �                    ECS|EPT|CamExtEnable   Enabled|Disabled   KEnables the cam signal to be extended by a specified number of crank pulses �     !              ECS|EPT|CamExtension   pulses   <Specifies the number of crank pulses to extend the cam pulse �                      ECS|EPT|CamHistory   #Normal|Error|Always High|Always Low   Cam Signal Status �                        ECS|EPT|CamOffset   pulses   <Specifies the number of crank pulses to offset the cam pulse �                      ECS|EPT|CamOffsetEnable   Enabled|Disabled   IEnables the cam signal to be offset by a specified number of crank pulses �     !              ECS|EPT|CamSelect   	Cam1|Cam2   (Selects which Cam signal is used for EPT �     !             ECS|EPT|CrankCount   pulses   #EPT crank pulse count while in sync �                        ECS|EPT|CrankRunThreshold   RPM   2Engine speed which determines EngineStatus=RUNNING �     	    C�            ECS|EPT|CrankStalled   |   *Indicates engine speed is below StallSpeed �     !              ECS|EPT|CrankSyncStopped   |   (Indicates EPT is not in sync with engine �     !              ECS|EPT|Crank_DigChanAsn_Mem       -Assigns digital signal source to crank signal �                    ECS|EPT|DI1-1_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                       ECS|EPT|DI1-2_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|DI2-1_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|DI2-2_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|DI3-1_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|DI3-2_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|DI4-1_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|DI4-2_TDC   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                      ECS|EPT|Dig_InvertConfig   usec   OSelects whether digital input is inverted before directed to channel assignment �                       ECS|EPT|Digital_Filt_Array   us   .Maximum time of rejected digital signal glitch �     	   @ ����       
                                               	   ECS|EPT|EPT_Type   "ENC Extrap 2|ENC Extrap 4|N-M |N+1   EPT Pattern Type Selection �                      ECS|EPT|EncZMask   EncZ Masked|EncZ Passed   lSelects whether encoder Z signal is masked by the selected cam signal or passed directly to the EPT function �     !             ECS|EPT|EngineSimEnable   |   %Enables simulation of select EPT type �     !              ECS|EPT|EngineSpeed   RPM   Indicates engine speed �     	                   ECS|EPT|EngineStatus   STALLED|CRANKING|RUNNING   7Engine status based on StallSpeed and CrankRunThreshold �                        ECS|EPT|GlobalTDCOffset   CAD   -Global TDC offset between absolute 0 and TDC1 �     	                  ECS|EPT|MaxCAT   CAT   3Maximum crank angle ticks for complete engine cycle �           �           ECS|EPT|MissedCamFlag   |   BIndicates that the EncZ rising edge was not detected when expected �     !               ECS|EPT|MissedCrankFlag   |   NIndicates that not enough crank pulses were received for complete engine cycle �     !               ECS|EPT|MissedGapFlag   |   ;Indicates that the crank gap was not detected when expected �     !               ECS|EPT|MissedPlus1Flag   |   CIndicates that the crank Plus1 pulse was not detected when expected �     !               ECS|EPT|NumberOfCrankTeeth   pulses   #Number of crank pulses per rotation �            <          ECS|EPT|NumberOfMissingTeeth   pulses   <Number missing adjacent crank teeth for the gap. M = 1 or 2. �                      ECS|EPT|Plus1Location   Retard|Advance   .Plus1 tooth location with respect to mid-point �     !             ECS|EPT|SimulatedSpeed   RPM   -Simulated engine speed during Simulation mode �     	    D            ECS|EPT|StallSpeed   RPM   BEngine speed at which EPT will lose sync and indicate CrankStalled �     	    A�            ECS|EPT|Stroke   4-STROKE|2-STROKE   Indicates 2 or 4-Stroke Engine �     !             ECS|EPT|SyncEnable   |   Enables EPT to sync �     !              ECS|EPT|SyncFlagClear   |   Clears EPT errors �     !              ECS|EPT|TDC1   CAD   Top Dead Center �     	                  ECS|EPT|TDC2   CAD   Top Dead Center �     	    Cp           ECS|EPT|TDC3   CAD   Top Dead Center �     	    C�           ECS|EPT|TDC4   CAD   Top Dead Center �     	    Bp           ECS|EPT|TDC5   CAD   Top Dead Center �     	    C�            ECS|EPT|TDC6   CAD   Top Dead Center �     	    D            ECS|EPT|TDC7   CAD   Top Dead Center �     	    B�           ECS|EPT|TDC8   CAD   Top Dead Center �     	    C�           ECS|Exec|CalVIEWInitOK   Failed|Success   1Indicates FPGA did not load.  Recompile required. �     !              ECS|Exec|Control_Duration   usec   Pulse generation process time �           �           ECS|Exec|MainLoopDuration   usec   Main RT loop execution time �           �           ECS|Exec|MainLoopPeriod   usec   Main RT loop period �           '           ECS|Exec|MainLoopPeriod_Set   usec   Main RT loop period setpoint �           '          ECS|Exec|Read_Inputs_Duration   usec   Pulse generation process time �           5            ECS|Exec|SlowSpeedLoopPeriod_Set   ms     �           �          ECS|Exec|Write_Outputs_Duration   usec   Pulse generation process time �           '           ECS|Faults|12V_Max       Maximum Voltage �     	                  ECS|Faults|12V_Min       Minimum Voltage �     	                  ECS|Faults|5V_Max       Maximum Voltage �     	                  ECS|Faults|5V_Min       Minimum Voltage �     	                  ECS|Faults|ECT_Max       Maximum Voltage �     	                  ECS|Faults|ECT_Min       Minimum Voltage �     	                  ECS|Faults|IAT_Max       Maximum Voltage �     	                  ECS|Faults|IAT_Min       Minimum Voltage �     	                  ECS|Faults|MAF_Max       Maximum Voltage �     	                  ECS|Faults|MAF_Min       Minimum Voltage �     	                  ECS|Faults|MAP_Max       Maximum Voltage �     	                  ECS|Faults|MAP_Min       Minimum Voltage �     	                  ECS|Faults|OilP_Max       Maximum Voltage �     	                  ECS|Faults|OilP_Min       Minimum Voltage �     	                  ECS|Faults|OilTemp_Max       Maximum Voltage �     	                  ECS|Faults|OilTemp_Min       Minimum Voltage �     	                  ECS|Faults|RPM_Max       Minimum Voltage �     	                  ECS|Faults|RailP_Max       Maximum Voltage �     	                  ECS|Faults|RailP_Min       Minimum Voltage �     	                  ECS|Faults|TDKBattV_Max       Maximum Voltage �     	                  ECS|Faults|TDKBattV_Min       Minimum Voltage �     	                  ECS|Fuel|AFStoich       %Air/Fuel mass ratio for stoichiometry �     	    Ak33           ECS|Fuel|AirDistributionArrayMAF   %   EMass air flow distribution for individual cylinders (must total 100%) �     	   @ ����                                                              	   ECS|Fuel|AirDistributionArraySD   %   ISpeed/Density air distribution for individual cylinders (must total 100%) �     	   @ ����                                              	   ECS|Fuel|AirMassArray   mg   !Air mass for individual cylinders �     	   @ ����                                                              	    ECS|Fuel|AirMassMAF   mg   MAF-based total air mass �     	                   ECS|Fuel|AirMassMode   MAF|SPEED/DENSITY   !Selects air mass calculation mode �                      ECS|Fuel|AirMassSD   mg   CSpeed-Density-based total theoretical air mass before Ve correction �     	                   ECS|Fuel|AirMassSDCorr   mg   6Speed-Density-based total air mass after Ve correction �     	                   ECS|Fuel|CalcAirDensity   Kg/m3   Air density �     	                   ECS|Fuel|ClosedLoopDieselFuel   Enabled|Disabled   2Enable closed loop control for the fuel quantities �     !              ECS|Fuel|CombustionMode   Diesel|Gasoline|Dual Fuel   Mode of Combustion Selection �                      ECS|Fuel|CrankingFuelEnrich   %/100   4Enrichment for fuel when engine is in cranking state �     	    ?��          ECS|Fuel|Cylinders       Number of cylinders �                     ECS|Fuel|DesDieselLambdaSetpoint       .Desired lambda setpoint before manual settings �     	                   ECS|Fuel|DesMainQuantity   mg   Desired main Quantity �     	                   ECS|Fuel|DesMainSOI   DBTDC   6Desired main start of injection before manual settings �     	                   ECS|Fuel|DesPilot1Quantity   mg   6Desired main start of injection before manual settings �     	                   ECS|Fuel|DesPilot1SOI   DBTDC   6Desired main start of injection before manual settings �     	    Bp             ECS|Fuel|DesPilot2Quantity   mg   6Desired main start of injection before manual settings �     	                   ECS|Fuel|DesPilot2SOI   DBTDC   6Desired main start of injection before manual settings �     	    Bp             ECS|Fuel|DesPost1Quantity   mg   6Desired main start of injection before manual settings �     	                   ECS|Fuel|DesPost1SOI   DBTDC   6Desired main start of injection before manual settings �     	    �p             ECS|Fuel|DesPost2Quantity   mg   6Desired main start of injection before manual settings �     	                   ECS|Fuel|DesPost2SOI   DBTDC   6Desired main start of injection before manual settings �     	    �p             ECS|Fuel|DieselFuelPIDOutput       4PID controller output (before feed forward is added) �     	                   ECS|Fuel|DieselLambdaSetpoint       -Final Labmda Setpoint used by the PID Control �     	                   ECS|Fuel|DieselLambdaTable   mm3/cyc|rpm|   Lambda setpoint lookup table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��       @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @   @             #ECS|Fuel|DieselManualLambdaSetpoint       Manual Lambda Setpoint �     	    @             )ECS|Fuel|DieselManualLambdaSetpointEnable   Enabled|Disabled   Enable Manual Lambda Setpoint �     !              ECS|Fuel|DieselPIDKp       Fuel PID Kp �     	                  ECS|Fuel|DieselPIDTd   min   Fuel PID Td �     	                  ECS|Fuel|DieselPIDTi   min   Fuel PID Ti �     	                  ECS|Fuel|ECTEnrichFactor       ECT enrichment factor �     	    >���           ECS|Fuel|ECTEnrichTable   C|   +Engine coolant temperature enrichment table �     	  @@ ����  X @@ ����  Y 
 P            A   A�  B   Bp  B�  B�  B�     >���>�ff?   ?L��?�  ?�  ?�  ?�            ECS|Fuel|EngineDisplacement   cc   Total engine displacement �     	    D�            ECS|Fuel|FuelMassCorr   mg   (Mass of Fuel injected per cylinder event �     	   @ ����                                                              	    ECS|Fuel|FuelPulseWidth   msec   !Final calculated fuel pulse width �     	   @ ����       @�  @�  @�  @�  @�  @�  @�  @�                         	    ECS|Fuel|FuelPulseWidthLimit   msec   Maximum permissable fuel pulse �     	    A             ECS|Fuel|InjCalibrationTable   mm3/inj|bar|usec   Fuel Injector Calibration �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             >L��?�  ?�  @   @   @@  @`  @�  @�  @�  @�  A   A   Ap  A�  A�  B   Bp  B�     BH  B�  B�  CH  Cz  C�  C�  D  DH  Dz  D�  D�� D�  D�� D�  D�  D�  D�@ D�` D�                                                                                               C� C�� C�  C�  C�  Cw  Cr  C}  Cz  Cx  Cv  Cu  Ct  Cf  Cf  Cf  Cf  Cf          D� C� C�  C�  C�  C�  C�  C�� C�  C�  C�  C�� C�  C{  C{  C{  C{  C{          D*� D  C� C�  C�� C�� C�� C�  C�� C�� C�� C�  C�� C�� C�� C�� C�� C��         D:@ D� D� C� C�  C�  C�� C�  C�� C�� C�� C�  C�� C�  C�  C�  C�  C�          DG@ D  D
� C�  C�  C�  C�� C�� C�  C�  C�  C�  C�  C�� C�� C�� C�� C��         DT� D%@ D  D  C� C�� C�� C�� C�  C�  C�  C�� C�� C�  C�  C�  C�  C�          Db  D/� D@ D� C� C C�� C�� C�  C�� C�  C�  C�� C�� C�� C�� C�� C��         Do@ D:@ D&� D  C�� C�  C�� C�� C�  C�� C�  C�� C�� C�� C�� C�� C�� C��         D�� DL� D7@ D'@ D� Cۀ CÀ C�� C�  C�� C�  C�� C�� C�  C�  C�  C�  C�          D�� D[  DC� D2� D� C�  Cр C�  C�� C�� C�� C�� C�� C�� C�� C�� C�� C��         D�` Dh� DO� D=� D  C�  C݀ Cƀ C�� C�� C�� C�  C�� C�  C�� C�� C�� C��         D�� Ds� DZ  DG  D � D  C�  C�  Cǀ C�  C�� C�  C�  C�  C�  C�  C�  C�          D�� D�` Dk  DV� D-� D@ C�  C�  C�  CӀ C�  C�  Cŀ C�  C�  C�  C�  C�          D�@ D�  D�� D{� DL  D � D� D  C�� C�  C� C�  Cۀ C�  C�  C�  C�  C�          D�� D�� D�  D�` Dg@ D7@ D  D@ D@ D� C�� C�  C� C� C� C� C� C�         E� D�@ D�@ D�` D�  D`@ D@� D-� D"  D@ D  D  D@ D  D  D  D  D          E&0 EP D�@ D�  D�  D�� Dc@ DJ  D:� D3� D-� D(� D#� D� D� D� D� D�         E;� E*� E� E` D�` D�� D�  D�� Do� De  D]  DU� DN� DC� DC� DC� DC� DC�         E;� E;� E;� E-0 E� D�` D�` D�� D�  D�� D�@ D�` D|@ Dm  Dm  Dm  Dm  Dm            ECS|Fuel|Inj_Pls_Switch       &Toggles ON/OFF each DI injection pulse �                    ECS|Fuel|InjectorOpen   msec   3Time for injector to open at current batery voltage �     	    @Mp�            ECS|Fuel|InjectorTurnOnTimeCoeff       /Coefficient for modifying injector turn on time �     	    ?(��          ECS|Fuel|LambdaCorr   Lambda   Corrected Lambda for bank 1 �     	    ?�             ECS|Fuel|LambdaPIDOut   Lambda    Lambda PID adjustment for bank 1 �     	                   ECS|Fuel|LambdaPID_Kc   Lambda/Lambda    Lambda control proportional gain �     	                  ECS|Fuel|LambdaPID_Max   Lambda   Maximum lambda PID adjustment �     	    >L��          ECS|Fuel|LambdaPID_Min   Lambda   Minimum lambda PID adjustment �     	    �L��          ECS|Fuel|LambdaPID_Td   min   Lambda control derivative time �     	                  ECS|Fuel|LambdaPID_Ti   min   Lambda control integral time �     	                  ECS|Fuel|LambdaTable   Kg/Hr|RPM|Lambda   Lambda Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             A�  B   Bp  B�  B�         Dz  D�  E;� Ez  E�@ E��       ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�  ?�            ECS|Fuel|LambdaTableOverride   MANUAL|TABLE   6TRUE uses ManualLambdaSetpoint; FALSE uses LambdaTable �     !              ECS|Fuel|MainQuantityTable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|MainSOITable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Man_FuelPulseWidth   msec   "fuel pulse width manual duty cycle �     	   @ ����       @�  @�  @�  @�  @�  @�  @�  @�                         	   ECS|Fuel|Man_PulseWidthOverride   |   Number of cylinders �     !             ECS|Fuel|ManualLambdaSetpoint   Lambda   +Manual setpoint for overriding lambda table �     	    ?�            ECS|Fuel|ManualMainDuration   DBTDC   Manual Main Start of Injection �     	    ?�            !ECS|Fuel|ManualMainDurationEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualMainSOI   DBTDC   Manual Main Start of Injection �     	                  ECS|Fuel|ManualMainSOIEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPFIFuelTiming   DBTDC   Manual fuel timing setpoint �     	                  ECS|Fuel|ManualPilot1Duration   msec   Manual Pilot Duration �     	                  #ECS|Fuel|ManualPilot1DurationEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPilot1SOI   DBTDC   Manual Main Start of Injection �     	    Bp            ECS|Fuel|ManualPilot1SOIEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPilot2Duration   msec   Manual Pilot 2 Duration �     	                  #ECS|Fuel|ManualPilot2DurationEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPilot2SOI   DBTDC   Manual Main Start of Injection �     	    Bp            ECS|Fuel|ManualPilot2SOIEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPost1Duration   msec    Manual Post 1 Injection Duration �     	                  "ECS|Fuel|ManualPost1DurationEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPost1SOI   DBTDC   Manual Main Start of Injection �     	    �             ECS|Fuel|ManualPost1SOIEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPost2Duration   msec   Manual Main Start of Injection �     	                  "ECS|Fuel|ManualPost2DurationEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|ManualPost2SOI   DBTDC   Manual Main Start of Injection �     	    �             ECS|Fuel|ManualPost2SOIEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !             ECS|Fuel|MaxTotalDieselFuel   mm3/cyc/cyl   Max Fuel Duty Cycle �     	                  ECS|Fuel|MinTotalDieselFuel   mm3/cyc/cyl   Min Fuel Duty Cycle �     	                  #ECS|Fuel|NextCycleFdBkControlEnable   Enabled|Disabled   %Enable Manual Main Start of Injection �     !              ECS|Fuel|PFIFuelControlMode   OPEN LOOP|WIDE BAND LAMBDA PID   Selects fuel control mode �                       ECS|Fuel|PFIFuelDensity   mg/cc   (Density of fuel at operating temperature �     	    D8N          ECS|Fuel|PFIFuelTiming   DBTDC   Final calculated fuel timing �     	    C             ECS|Fuel|PFIFuelTimingTable_MAF   Kg/Hr|RPM|DBTDC   (Fuel Timing Table based on Speed and MAF �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             CH  C�  D  DH  Dz         Dz  D�  E;� Ez  E�@ E��       C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C            ECS|Fuel|PFIFuelTimingTable_MAP   kPa|RPM|DBTDC   (Fuel Timing Table based on Speed and MAP �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             CH  C�  D  DH  Dz         Dz  D�  E;� Ez  E�@ E��       C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C  C            ECS|Fuel|PFIInjectorFlowRate   cc/min   Nominal injector flow rate �     	    CM            ECS|Fuel|PFIInjectorOpenTable   V|msec   Injector opening time table �     	  @@ ����  X @@ ����  Y 
 P        @�  @�  A   A  A   A0  A@  AP  A`  Ap  A�     @Mp�@*=q@��?��H?�(�?��
?���?�  ?��?�ff?xQ�          ECS|Fuel|PFITableFuelTiming   |   3F = Use FuelTimingSetpoint; T = Use TableFuelTiming �     !             ECS|Fuel|PID_FuelPulseWidth   msec   !Final calculated fuel pulse width �     	   @ ����       @�%@�%@�%@�%@�%@�%@�%@�%@�%@�%@�%@�%       	    ECS|Fuel|Pilot1QuantityTable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Pilot1SOITable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Pilot2QuantityTable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A�            ECS|Fuel|Pilot2SOITable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Post1QuantityTable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Post1SOITable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Post2QuantityTable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|Post2SOITable   mm3/cyc|rpm|DBTDC   $Main Start of Injection Lookup Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E;� EZ� Ej` Ez  E�� E��               �� ��     ?� @  @ �@@  @_�
@�?�A/�A\�A�  A���A��        �� �� �� T>� T>� T>� T?���?�  @@  A/�A\�A�  A��A��        ����� ����    >� T?���?���?�  @@  A/�A\�A�  A��A��        ������ T�� T    >� T?���?�  ?� @`��A/�A\�A�  A��A��                    >� T?���?�  ?�  ?� @`��A/�A\�A�  A��A���    >���>� T>� T>� T?���?�  ?�  ?� ?� @`��A/�A\�A�  A��A��    >� T?���?���?���?���?�  ?�  ?� ?� @�?�A4  A\�A�  A��A���    ?@  ?���?���?���?���?� ?� ?� @ �@�?�A8�A_�A�  A��A��    ?���?�  ?�  ?�  ?�  ?� @ �@ �@@  @�?�A;�Ad  A���A���A���?���?� ?� ?� ?� ?� @ �@@  @@  @_�
@��AF  Ah�A���A�� A���?���?� @ �@ �@ �@ �@@  @_�
@�?�@�  @�?�AP�Ax��A�0A���A�O�?���?� @/�
@_�
@@  @@  @�?�@�?�@�  @�  A  Ae�A���A�@ A���A�� ?���?� @/�
@_�
@_�
@�?�@�  @��@�  @�?�A(  Am��A��A��A�@ A��?���?� @/�
@_�
@�  @�?�@�?�@�  @�  A�A8�Aw�A���A�  A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��?���?� @/�
@_�
@�  @�?�@�?�@��A�A�AG�A��A��A��A��A��          ECS|Fuel|VeTable   	kPa|RPM|%   Volumetric Efficiency Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             A�  B   Bp  B�  B�         Dz  D�  E;� Ez  E�@ E��       B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�  B�            ECS|Inputs|12VPulsBattV   V   12V Supply Voltage �     	    <��           ECS|Inputs|5VPulsBattV   V   5V Supply Voltage �     	    >�@           ECS|Inputs|Coolant_Temp       *Coolant temperature from calibration table �     	                   ECS|Inputs|Coolant_Temp_Conv   V|%   %Coolant temperature calibration table �     	  @@ ����  X @@ ����  Y 
 P            @�         B�            #ECS|Inputs|Coolant_Temp_FilterBreak   Hz   +Coolant temperature filter cutoff frequency �     	    A�            ECS|Inputs|Coolant_Temp_Raw       Raw coolant temperature reading �     	    �zN=           ECS|Inputs|ECT       ECT from calibration table �     	                   ECS|Inputs|ECT_Conv   V|%   ECT calibration table �     	  @@ ����  X @@ ����  Y 
 P            @�         B�            ECS|Inputs|ECT_FilterBreak   Hz   ECT filter cutoff frequency �     	    A�            ECS|Inputs|ECT_Raw       Raw ECT reading �     	    �zN=           ECS|Inputs|EGR1_Pos       $EGR1 Position from calibration table �     	    ?              ECS|Inputs|EGR1_Pos_Conv   V|   EGR1 Position Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            ECS|Inputs|EGR1_Pos_FilterBreak   Hz   %EGR1 Position Filter cutoff frequency �     	    A�            ECS|Inputs|EGR1_Pos_Raw       Output from calibration table �     	    <�             ECS|Inputs|EGRc_P_in       Output from calibration table �     	    ?              ECS|Inputs|EGRc_P_in_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�             ECS|Inputs|EGRc_P_in_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|EGRc_P_in_Raw       Output from calibration table �     	    <�             ECS|Inputs|EGRc_P_out       Output from calibration table �     	    ?              ECS|Inputs|EGRc_P_out_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            !ECS|Inputs|EGRc_P_out_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|EGRc_P_out_Raw       Output from calibration table �     	    <�             #ECS|Inputs|Enable_Coolant_Temp_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_ECT_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_EGR1_Pos_Filt   Enable|Disable   Enable use of filter �     !               ECS|Inputs|Enable_EGRc_P_in_Filt   Enable|Disable   Enable use of filter �     !              !ECS|Inputs|Enable_EGRc_P_out_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_IAT_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_MAF_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_MAP_Filt   Enable|Disable   Enable use of filter �     !               ECS|Inputs|Enable_Oil_Press_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_Oil_Temp_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_Pedal_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|Enable_RailP_Filt   Enable|Disable   Enable use of filter �     !              !ECS|Inputs|Enable_Turbo_P_in_Filt   Enable|Disable   Enable use of filter �     !              "ECS|Inputs|Enable_Turbo_P_out_Filt   Enable|Disable   Enable use of filter �     !              ECS|Inputs|IAT       Output from calibration table �     	                   ECS|Inputs|IAT_Conv   V|%   Calibration table �     	  @@ ����  X @@ ����  Y 
 P            @�         B�            ECS|Inputs|IAT_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|IAT_Raw       Output from calibration table �     	    �zN`           !ECS|Inputs|Init_Coolant_Temp_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_ECT_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_EGR1_Pos_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_EGRc_P_in_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_EGRc_P_out_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_IAT_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_MAF_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_MAP_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_Oil_Press_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_Oil_Temp_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_Pedal_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_RailP_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|Init_Turbo_P_in_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !               ECS|Inputs|Init_Turbo_P_out_Filt   Enable|Disable   -Re-intialize filter to change break frequency �     !              ECS|Inputs|MAF       Output from calibration table �     	    ?              ECS|Inputs|MAF_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            ECS|Inputs|MAF_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|MAF_Raw       Output from calibration table �     	    =/             ECS|Inputs|MAP       Output from calibration table �     	    ?              ECS|Inputs|MAP_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            ECS|Inputs|MAP_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|MAP_Raw       Output from calibration table �     	    <�             ECS|Inputs|Oil_Press       Output from calibration table �     	    ?              ECS|Inputs|Oil_Press_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�             ECS|Inputs|Oil_Press_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|Oil_Press_Raw       Output from calibration table �     	    <�             ECS|Inputs|Oil_Temp       Output from calibration table �     	                   ECS|Inputs|Oil_Temp_Conv   V|%   Calibration table �     	  @@ ����  X @@ ����  Y 
 P            @�         B�            ECS|Inputs|Oil_Temp_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|Oil_Temp_Raw       Output from calibration table �     	    �zN=           ECS|Inputs|Pedal       Output from calibration table �     	    A���           ECS|Inputs|Pedal_Conv   V|%   Calibration table �     	  @@ ����  X @@ ����  Y 
 P            @�         B�            ECS|Inputs|Pedal_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|Pedal_Raw       Output from calibration table �     	    <�             ECS|Inputs|RailP       Output from calibration table �     	    ?              ECS|Inputs|RailP_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            ECS|Inputs|RailP_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|RailP_Raw       Output from calibration table �     	    <�             !ECS|Inputs|SimEnable_Coolant_Temp   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_ECT   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_EGR1_Pos   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_EGRc_P_in   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_EGRc_P_out   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_IAT   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_MAF   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_MAP   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_Oil_Press   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_Oil_Temp   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_Pedal   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !             ECS|Inputs|SimEnable_RailP   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|SimEnable_Turbo_P_in   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !               ECS|Inputs|SimEnable_Turbo_P_out   Enabled|Disabled   8Enable simulation of this parameter in engineering units �     !              ECS|Inputs|Sim_Coolant_Temp       Simulation value �     	                  ECS|Inputs|Sim_ECT       Simulation value �     	                  ECS|Inputs|Sim_EGR1_Pos       Simulation value �     	                  ECS|Inputs|Sim_EGRc_P_in       Simulation value �     	                  ECS|Inputs|Sim_EGRc_P_out       Simulation value �     	                  ECS|Inputs|Sim_IAT       Simulation value �     	                  ECS|Inputs|Sim_MAF       Simulation value �     	                  ECS|Inputs|Sim_MAP       Simulation value �     	                  ECS|Inputs|Sim_Oil_Press       Simulation value �     	                  ECS|Inputs|Sim_Oil_Temp       Simulation value �     	                  ECS|Inputs|Sim_Pedal       Simulation value �     	    A���          ECS|Inputs|Sim_RailP       Simulation value �     	                  ECS|Inputs|Sim_Turbo_P_in       Simulation value �     	                  ECS|Inputs|Sim_Turbo_P_out       Simulation value �     	                  ECS|Inputs|TDKBattV   V   TDK Battery Voltage �     	    =hw           ECS|Inputs|Turbo_P_in       Output from calibration table �     	    ?              ECS|Inputs|Turbo_P_in_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            !ECS|Inputs|Turbo_P_in_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|Turbo_P_in_Raw       Output from calibration table �     	    <�             ECS|Inputs|Turbo_P_out       Output from calibration table �     	    ?              ECS|Inputs|Turbo_P_out_Conv   V|   Calibration table �     	  @@ ����  X @@ ����  Y 
 P        ?   @�     ?   @�            "ECS|Inputs|Turbo_P_out_FilterBreak   Hz   Filter cutoff frequency �     	    A�            ECS|Inputs|Turbo_P_out_Raw       Output from calibration table �     	    <�             ECS|MAF|DesHP-EGR%Open   %   ,Desired EGR Duty Cycle before Manual Setting �     	    B�             ECS|MAF|DesMAF   Kg/Hr   *Desired MAF Setpoint before Manual Setting �     	    BX             ECS|MAF|HP-EGRDC   %   Final Boost Duty Cycle �     	                   ECS|MAF|HP-EGRDCTable   %|%Open   EGR Duty Cycle Map �     	  @@ ����  X @@ ����  Y 
 P        <G�=��B��B�     B�  B�  @�  @�            ECS|MAF|LP-EGRDC   %   Final Boost Duty Cycle �     	                   ECS|MAF|MAFBaseDesTable   mm3/cyc|rpm|Kg/Hr   Base MAF Setpoint Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B  B  B   B*     D;� DR  Dz  D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ� E��       BX  A��TB��B7  B[��BoffB�33B���C  C� C%��C�  C�  D  BX  A��#BffB4  BP��B^��B�  B���C  CL�C"  C�  C�  D  BX  A��#B��B(  BX  BZffBy��B�ffB�  C �3C��C�  C�  D  Ba  A��B  B4  BX  BoffB�ffB�  B�  CL�C%��C�  C�  D  Bs  B&�B(  B:  B_33B�33B�ffB�  B�  C33C.��C�  C�  D  B���B/dZB;33BR  Bq33B��3B���Bҙ�C  C�C;33C�  C�  D  B�� BO��BS33Bg  B���B�33B�  B���C� C%  CG��C�  C�  D  B��fBk�;Bk33B�� B���B��B�  B���C  C+��CO  C�  C�  D  B�  B�{B�  B�  B���B�33B홚CY�C"  C7&fC[��C�  C�  D  B�  B�;dB�
=B�  B�33B�ffB�ffC��C)� CA�Cj  C�  C�  D  B�  B�l�B�  Bʀ B���B�C33C��C1  CG�fCxffC�  C�  D  B�  Bϥ�B���B� B���CL�C  C#Y�C@  CY��C���C�  C�  D  B�  B��
B�  C� B���C�C ��C3��CR  Ct33C�� C�  C�  D  B�  B��TC
��C  C��C*�C1��CG��Cg  C���C�33C�  C�  D  B�  B��C33C� C;33C\� C�ffC��fC�@ C��fC���C�  C�  D  B�  B��C  C4  CX  C|  C�  C�  C�  C�  C�  C�  C�  D            ECS|MAF|MAFControlKp       
MAF PID Kp �     	                  ECS|MAF|MAFControlTd   min   
MAF PID Td �     	                  ECS|MAF|MAFControlTi   min   
MAF PID Ti �     	                  ECS|MAF|MAFCorrEnable   Corrected|Not Corrected   Enables MAF Correction �     !              ECS|MAF|MAFCorrTable   mm3/cyc|rpm|mg/cyl   MAF Correction Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B  B  B   B*     D;� DR  Dz  D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ� E��       D/  D/  D/  DC  DR  D\  Df  D�� D�  D�@ D�@ D�@ D�@ D�@ D/  D/  D/  DE� DT� D^� Df  D�� D�  D�@ D�@ D�@ D�@ D�@ D/  D/  D/  DE� DW  D^� Df  D�� D�  D�@ D�@ D�@ D�@ D�@ D/  D/  D/  DE� DY� D^� Dh� D�� D�  D�@ D�@ D�@ D�@ D�@ D/  D/  D/  DH  D\  Dc� Dm� D�� D�  D�@ D�@ D�@ D�@ D�@ D1� D1� D1� DJ� Da  Dp  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Df  D�� D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@ D4  D4  D4  DM  Dh� D�  D�� D�� D�  D�@ D�@ D�@ D�@ D�@           ECS|MAF|MAFECTCorrTable   C|   !MAF correction table based on ECT �     	  @@ ����  X @@ ����  Y 
 P        
��  �       Ap  A�  B  B4  B\  B�  B�     
?�  ?�  ?�  >��=�\)=u=#�
<��
                  ECS|MAF|MAFPIDEnable   |   Enable MAF PID �     !              ECS|MAF|MAFSetpoint   Kg/Hr   MAF PID Setpoint �     	    BX             ECS|MAF|ManualHP-EGR%DC   %   Manual EGR Duty Cycle Setting �     	                  ECS|MAF|ManualHP-EGREnable   Manual|Automatic   +Override EGR duty cycle with manual setting �     !             ECS|MAF|ManualLP-EGRDC   %   Manual EGR Duty Cycle Setting �     	                  ECS|MAF|ManualMAFSetpoint   Kg/Hr   Manual MAF Setting �     	                  ECS|MAF|ManualMAFSetpointEnable   Manual|Automatic   )Override MAF setpoint with manual setting �     !              ECS|MAF|MaxHP-EGR%DC    %   Max EGR Opening �     	                  ECS|MAF|MaxLP-EGRDC   %   Max EGR Opening �     	                  ECS|MAF|Max_PID_HP-EGRDC   %   Max EGR Opening �     	                  ECS|MAF|MinHP-EGR%DC   %   Min EGROpening �     	                  ECS|MAF|MinLP-EGRDC   %   Min EGROpening �     	                  ECS|MAF|Min_PID_HP-EGRDC   %   Min EGROpening �     	                  ECS|NextCycle|MFBPIDKc   DBTDC   Spark Operating Window Start �     	                  ECS|NextCycle|MFBPIDOutputHigh   DBTDC   Spark Operating Window Start �     	                  ECS|NextCycle|MFBPIDOutputLow   DBTDC   Spark Operating Window Start �     	                  ECS|NextCycle|MFBPIDTd   DBTDC   Spark Operating Window Start �     	                  ECS|NextCycle|MFBPIDTi   DBTDC   Spark Operating Window Start �     	                  ECS|NextCycle|MFBPIDTimeout   msec   &Timeout in msec for Next Cycle Control �            d          ECS|NonCriticalFault|DI1   Error|OK   Non Critical Fault �     !               ECS|NonCriticalFault|DI2   Error|OK   Non Critical Fault �     !               ECS|NonCriticalFault|DI3   Error|OK   Non Critical Fault �     !               ECS|NonCriticalFault|DI4   Error|OK   Non Critical Fault �     !               ECS|NonCriticalFault|PFI1   Error|OK   Non Critical Fault �     !               ECS|NonCriticalFault|PFI2   Error|OK   Non Critical Fault �     !               #ECS|NonCriticalFault|Throttle1Fault   Error|OK   Non Critical Fault �     !              ECS|NonCriticalFault|UEGO   Error|OK   Non Critical Fault �     !              ECS|NonCriticalFault|UEGO2   Error|OK   Non Critical Fault �     !              "ECS|PFI1|PFI1_LS1_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI1|PFI1_LS1_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               "ECS|PFI1|PFI1_LS2_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI1|PFI1_LS2_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               "ECS|PFI1|PFI1_LS3_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI1|PFI1_LS3_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               "ECS|PFI1|PFI1_LS4_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI1|PFI1_LS4_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               ECS|PFI1|PFI1_ModulePresent   ON|OFF   :Indicates PFI Driver module present and externally powered �     !               ECS|PFI1|PFI1_ModuleRev       0Indicates DI Driver module Hardware/Firmware Rev �     0����                  ECS|PFI1|PFI1_OpenFaultOverride   Override|Show Fault   4Determines whether open-circuit faults are indicated �     !              "ECS|PFI1|PFI1_PF11OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               "ECS|PFI1|PFI1_PF12OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               "ECS|PFI1|PFI1_PF13OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               "ECS|PFI1|PFI1_PF14OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               #ECS|PFI1|PFI1_PFI1ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               #ECS|PFI1|PFI1_PFI2ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               #ECS|PFI1|PFI1_PFI3ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               #ECS|PFI1|PFI1_PFI4ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               "ECS|PFI2|PFI2_LS1_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI2|PFI2_LS1_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               "ECS|PFI2|PFI2_LS2_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI2|PFI2_LS2_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               "ECS|PFI2|PFI2_LS3_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI2|PFI2_LS3_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               "ECS|PFI2|PFI2_LS4_OpenCircuitFault   ON|OFF   "Lowside channel open-circuit fault �     !               #ECS|PFI2|PFI2_LS4_ShortCircuitFault   ON|OFF   #Lowside channel short-circuit fault �     !               ECS|PFI2|PFI2_ModulePresent   ON|OFF   :Indicates PFI Driver module present and externally powered �     !               ECS|PFI2|PFI2_ModuleRev       0Indicates DI Driver module Hardware/Firmware Rev �     0����                  ECS|PFI2|PFI2_OpenFaultOverride   Override|Show Fault   4Determines whether open-circuit faults are indicated �     !              "ECS|PFI2|PFI2_PF11OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               "ECS|PFI2|PFI2_PF12OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               "ECS|PFI2|PFI2_PF13OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               "ECS|PFI2|PFI2_PF14OpenCircuitFault   ON|OFF   Injector open-circuit fault �     !               #ECS|PFI2|PFI2_PFI1ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               #ECS|PFI2|PFI2_PFI2ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               #ECS|PFI2|PFI2_PFI3ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               #ECS|PFI2|PFI2_PFI4ShortCircuitFault   ON|OFF   Injector short-circuit fault �     !               ECS|PFI|I_Duration   msec   Duration for this phase �     	   @ ����       ?�      ?�      ?�      ?�             	   ECS|PFI|I_Setpoint   A   Current setpoint for this phase �     	   @ ����       @@  ?�  @@  ?�  @@  ?�  @@  ?�         	   ECS|PFI|PFICutOffPosition   CAD   -Global TDC offset between absolute 0 and TDC1 �     	    �p            ECS|PFI|PFIMod1_FaultClear   	Clear|OFF     �     !              ECS|PFI|PFIMod1_ModuleEnable   ON|OFF     �     !              ECS|PFI|PFIMod1_OneShot   ON|OFF     �     !              ECS|PFI|PFIMod1_OneShotDuration   msec     �     	    @�            ECS|PFI|PFIMod1_OneShotSelect   Disabled|PFI1|PFI2|PFI3|PFI4     �                      ECS|PFI|PFIMod1_PFI1_Enable   Enabled|Disabled     �     !             *ECS|PFI|PFIMod1_PFI1_Phase1FirstPeakEnable   ON|OFF     �     !             !ECS|PFI|PFIMod1_PFI1_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|PFI|PFIMod1_PFI2_Enable   Enabled|Disabled     �     !             *ECS|PFI|PFIMod1_PFI2_Phase1FirstPeakEnable   ON|OFF     �     !             !ECS|PFI|PFIMod1_PFI2_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|PFI|PFIMod1_PFI3_Enable   Enabled|Disabled     �     !             *ECS|PFI|PFIMod1_PFI3_Phase1FirstPeakEnable   ON|OFF     �     !             !ECS|PFI|PFIMod1_PFI3_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|PFI|PFIMod1_PFI4_Enable   Enabled|Disabled     �     !             *ECS|PFI|PFIMod1_PFI4_Phase1FirstPeakEnable   ON|OFF     �     !             !ECS|PFI|PFIMod1_PFI4_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|PFI|PFIMod2_FaultClear   	Clear|OFF     �     !              ECS|PFI|PFIMod2_ModuleEnable   ON|OFF     �     !              ECS|PFI|PFIMod2_OneShot   ON|OFF     �     !              ECS|PFI|PFIMod2_OneShotDuration   msec     �     	                  ECS|PFI|PFIMod2_OneShotSelect   Disabled|PFI1|PFI2|PFI3|PFI4     �                       ECS|PFI|PFIMod2_PFI1_Enable   Enabled|Disabled     �     !              *ECS|PFI|PFIMod2_PFI1_Phase1FirstPeakEnable   ON|OFF     �     !              !ECS|PFI|PFIMod2_PFI1_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|PFI|PFIMod2_PFI2_Enable   Enabled|Disabled     �     !              *ECS|PFI|PFIMod2_PFI2_Phase1FirstPeakEnable   ON|OFF     �     !              !ECS|PFI|PFIMod2_PFI2_RecircAlways   4-STROKE|2-STROKE     �     !              ECS|PFI|PFIMod2_PFI3_Enable   Enabled|Disabled     �     !              *ECS|PFI|PFIMod2_PFI3_Phase1FirstPeakEnable   4-STROKE|2-STROKE     �     !              !ECS|PFI|PFIMod2_PFI3_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|PFI|PFIMod2_PFI4_Enable   Enabled|Disabled     �     !              *ECS|PFI|PFIMod2_PFI4_Phase1FirstPeakEnable   ON|OFF     �     !              !ECS|PFI|PFIMod2_PFI4_RecircAlways   Recirc ON|Recirc OFF     �     !              ECS|RPC|BattV   V   0Battery voltage measured by the DI Driver module �     	    =hw           ECS|RPC|HPV_Current   A   QEstimated current to HPV based on battery voltage and nominal solenoid resistance �     	                   ECS|RPC|HPV_DC   %   Final HPV duty cycle �     	                   ECS|RPC|HPV_Enable   |   Enables PWM control of HPV �     !              ECS|RPC|HPV_Freq   Hz   &Operating Frequency of HPV PWM command �     	    Dz            ECS|RPC|HPV_Kc   %/bar   HPV PID proportional gain �     	    :�o          ECS|RPC|HPV_Kp_Action   %   /Proportional contribution of HPV PID controller �     	                   ECS|RPC|HPV_ManualDC   %   ?Value to override HPV PID final output when ManualOverride=TRUE �     	                  ECS|RPC|HPV_ManualOverride   |   0Causes ManualDC to override HPV PID final output �     !              ECS|RPC|HPV_MaxDC   %   XMaximum allowed duty cycle for HPV. This value is effective if lower than HPV_MaxDCCalc. �     	                  ECS|RPC|HPV_MaxDCCalc   %   �Maximum allowed duty cycle for HPV based on battery voltage and nominal solenoid resistance to limit current to 3A for channel pair �     	                   ECS|RPC|HPV_MinDC   %   "Minimum allowed duty cycle for HPV �     	                  ECS|RPC|HPV_NomResistance   Ohms   "Nominal resistance of HPV solenoid �     	    @@            ECS|RPC|HPV_NonPIDFF   %   FDuty cycle feed forward for the HPV while doing PID control of the IMV �     	    B             ECS|RPC|HPV_PID   %   pHPV PID controller output added to HPVPIDFF. Result is directed to selected PFI LS channel duty cycle parameter. �     	                   ECS|RPC|HPV_PIDFF   %   3Duty cycle feed forward added to the HPV PID output �     	    A�            ECS|RPC|HPV_PIDMax   %   ;HPV PID output maximum limit (before feed forward is added) �     	    A�            ECS|RPC|HPV_PIDMin   %   ;HPV PID output minimum limit (before feed forward is added) �     	    ��            ECS|RPC|HPV_Td   min   YDerivative time constant for HPV PID controller (higher = stronger action. 0 = disabled.) �     	                  ECS|RPC|HPV_Td_Action   A   -Derivative contribution of HPV PID controller �     	                   ECS|RPC|HPV_Ti   min   VIntegral time constant for HPV PID controller (lower = stronger action. 0 = disabled.) �     	                  ECS|RPC|HPV_Ti_Action   %   +Integral contribution of HPV PID controller �     	                   ECS|RPC|IMV_Current   A   QEstimated current to IMV based on battery voltage and nominal solenoid resistance �     	                   ECS|RPC|IMV_DC   %   Final IMV duty cycle �     	                   ECS|RPC|IMV_Enable   |   Enables PWM control of IMV �     !              ECS|RPC|IMV_Freq   Hz   &Operating Frequency of IMV PWM command �     	    C/            ECS|RPC|IMV_Kc   %/bar   IMV PID proportional gain �     	    :�o          ECS|RPC|IMV_Kp_Action   %   /Proportional contribution of IMV PID controller �     	                   ECS|RPC|IMV_ManualDC   %   ?Value to override IMV PID final output when ManualOverride=TRUE �     	                  ECS|RPC|IMV_ManualOverride   |   0Causes ManualDC to override IMV PID final output �     !              ECS|RPC|IMV_MaxDC   %   XMaximum allowed duty cycle for IMV. This value is effective if lower than IMV_MaxDCCalc. �     	                  ECS|RPC|IMV_MaxDCCalc   %   �Maximum allowed duty cycle for IMV based on battery voltage and nominal solenoid resistance to limit current to 3A for channel pair �     	                   ECS|RPC|IMV_MinDC   %   "Minimum allowed duty cycle for IMV �     	                  ECS|RPC|IMV_NomResistance   Ohms   "Nominal resistance of IMV solenoid �     	    @             ECS|RPC|IMV_NonPIDFF   %   FDuty cycle feed forward for the IMV while doing PID control of the HPV �     	    A�            ECS|RPC|IMV_PID   %   pIMV PID controller output added to IMVPIDFF. Result is directed to selected PFI LS channel duty cycle parameter. �     	                   ECS|RPC|IMV_PIDFF   %   3Duty cycle feed forward added to the IMV PID output �     	    A�            ECS|RPC|IMV_PIDMax   %   ;IMV PID output maximum limit (before feed forward is added) �     	    A�            ECS|RPC|IMV_PIDMin   %   ;IMV PID output minimum limit (before feed forward is added) �     	    ��            ECS|RPC|IMV_Td   min   YDerivative time constant for IMV PID controller (higher = stronger action. 0 = disabled.) �     	                  ECS|RPC|IMV_Td_Action   A   -Derivative contribution of IMV PID controller �     	                   ECS|RPC|IMV_Ti   min   VIntegral time constant for IMV PID controller (lower = stronger action. 0 = disabled.) �     	                  ECS|RPC|IMV_Ti_Action   %   +Integral contribution of IMV PID controller �     	                   "ECS|RPC|ManualEnableRailP_Setpoint   |   Enables PWM control of IMV �     !              ECS|RPC|Manual_RailP_Setpoint   bar   /Manual Rail pressure setpoint to PID controller �     	                  ECS|RPC|PFIBattV   (TDK 1U Rack Supply|12V Puls Power Supply   -Selects Power Supply Source for PFI/LS Module �                       ECS|RPC|RPC_FaultClear   #Clear RailP Fault|Clear RailP Fault   .Clears faults related to rail pressure control �     !              ECS|RPC|RailP   bar   Rail pressure in bar �     	    ?              ECS|RPC|RailP_ControlMode   IMV PID MODE|HPV PID MODE   +Selects the IMV or HPV as controlled by PID �                       ECS|RPC|RailP_Fault   Fault|No Fault   (Indicates the rail pressure fault status �     !               ECS|RPC|RailP_Max_Thresh   bar   hRail pressure maximum threshold which causes a critical fault and shuts down associated PFI LSX channels �     	    D�            ECS|RPC|RailP_Setpoint   bar   Final rail pressure Setpoint �     	    C�             ECS|RPC|RailP_Table   mm3/cyc|rpm|bar   $Injection Pressure calibration table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         @�  A   A   AP  Ap  A�  A�  A�  A�  A�  A�  B  B   BH  Bp  B�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ� Ez  E��       C�  C�  C�  C�  C�  Cπ C�  D@ D@ D  D@ D� D@ D� D!@ D!@ C�  C�  C�  C�  C�  C�  D	� D� D"� D'� D'� D'� D'� D'� D'� D(� C�  C�  C�  C�  C�  D	� D  D4  D9  D;� D;� D;� D;� D;� D;� D;� C�  C�  C�� C�  C�  D  D*  D@� DE� DH  DH  DH  DH  DH  DH  DH  C�  C�  C�� C�  C�  D"� D6� DM  DT� D\  D\  D\  D\  D\  D\  D\  C�  C�  C�  C�  D  D4  DJ� D\  Df  Dm� Dm� Dm� Dm� Dm� Dm� Dm� C�  C�  C�� C�  D  DC  D^� Dr� Dz  Dz  Dz  Dz  Dz  D|� D  D  C�  C�� C�  D  D  DH  Dc� Dw� D  D�� D�` D�  D�@ D�� D�  D�  C�  C�� CԀ D	� D%  DM  Dh� D|� D�  D�� D�� D�� D�� D�  D�� D�� C�  C�  Cހ D� D/  DR  Dm� D�� D�� D�� D�  D�� D�@ D�  D�� D�� C�  C�  C�  D  D@� DW  Dr� D�@ D�� D�� D�@ D�  D�  D�  D�� D�� C�  C�  C�  D/  DR  Da  Dz  D�  D�� D�  D�  D�� D�@ D�@ D�  D�@ C�  C�  C�  DC  Df  Dk  D�  D�@ D�� D�@ D�� D�  D�� D�� D�� D�  C�  C�  C�  DC  Df  D|� D�� D�� D�@ D�� D�@ D�� D�  D�  D�  D�  C�  C�  C�  DC  Df  D�  D�� D�� D�� D�@ D�� D�  D�  D�  D�  D�  C�  C�  C�  DC  Df  D�  D�� D�� D�� D�@ D�� D�  D�  D�  D�  D�            ECS|Scope|DI1_Scope       "DI Scope current and voltage trace �     	   @ ��������                     
    ECS|Scope|DI1_ScopeRefresh   REFRESH|OFF   Refreshes DI scope data �     !              ECS|Scope|DI2_Scope       "DI Scope current and voltage trace �     	   @ ��������                     
    ECS|Scope|DI2_ScopeRefresh   REFRESH|OFF   Refreshes DI scope data �     !              ECS|Scope|DI3_Scope       "DI Scope current and voltage trace �     	   @ ��������                     
    ECS|Scope|DI3_ScopeRefresh   REFRESH|OFF   Refreshes DI scope data �     !              ECS|Scope|DI4_Scope       "DI Scope current and voltage trace �     	   @ ��������                     
    ECS|Scope|DI4_ScopeRefresh   REFRESH|OFF   Refreshes DI scope data �     !              ECS|Sensors|UEGO Filter   Hz     �     	    ?�            ECS|Spark|Delay1   DBTDC   Spark Operating Window Start �     	    =���          ECS|Spark|Delay2   DBTDC   Spark Operating Window Start �     	    =���          ECS|Spark|Delay3   DBTDC   Spark Operating Window Start �     	    =���          ECS|Spark|MainMaxDwell   msec   Spark Operating Window Start �     	    A             ECS|Spark|MainSparkDwell   msec   Final calculated spark dwell �     	    @@             ECS|Spark|ManualSparkMainDwell   msec   Manual spark timing setpoint �     	    @@            ECS|Spark|ManualSparkTiming   DBTDC   Manual spark timing setpoint �     	                  ECS|Spark|Restrike1Dwell    msec   Spark Operating Window Start �     	    ?�            ECS|Spark|Restrike1Enable   |   Spark Operating Window Start �     !              ECS|Spark|Restrike2Dwell   msec   Spark Operating Window Start �     	    ?�            ECS|Spark|Restrike2Enable   |   Spark Operating Window Start �     !              ECS|Spark|Restrike3Dwell   msec   Spark Operating Window Start �     	    ?�            ECS|Spark|Restrike3Enable   |   Spark Operating Window Start �     !              ECS|Spark|RevLimitSparkRetard   CAD   -Degrees to retard when NCF rev limiter is hit �     	    A�            ECS|Spark|Spark1Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark2Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark3Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark4Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark5Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark6Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark7Enable   ON|OFF   Spark enable �     !              ECS|Spark|Spark8Enable   ON|OFF   Spark enable �     !              ECS|Spark|SparkDwellTable   V|msec   ,Spark dwell as a function of battery voltage �     	  @@ ����  X @@ ����  Y 
 P        @�  @�  A   A  A   A0  A@  AP  A`  Ap  A�     @�  @���@�33@���@�ff@�  @s33@fff@Y��@L��@@            ECS|Spark|SparkTiming   DBTDC   Final calculated spark timing �     	                   ECS|Spark|SparkTimingTable_MAF   Kg/Hr|RPM|DBTDC   )Spark Timing Table based on Speed and MAF �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             CH  C�  D  DH  Dz         Dz  D�  E;� Ez  E�@ E��       A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�            ECS|Spark|SparkTimingTable_MAP   kPa|RPM|DBTDC   )Spark Timing Table based on Speed and MAP �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             CH  C�  D  DH  Dz         Dz  D�  E;� Ez  E�@ E��       A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�  A�            ECS|Spark|Spark_Window_End   DBTDC   Spark Operating Window Start �     	    ´            ECS|Spark|Spark_Window_Start   DBTDC   Spark Operating Window Start �     	    B�            ECS|Spark|TableSparkMainDwell   Table|Manual   <F = Use SparkMainDwell Setpoint; T = Use TableSparkMainDwell �     !              ECS|Spark|TableSparkTiming   Table|Manual   5F = Use SparkTimingSetpoint; T = Use TableSparkTiming �     !              ECS|System|Power_Enable   |   &Enables DC all DC power to I/O drawers �     !              ECS|Throttle1|Chan1ControlMode   Position Feedback|Open Loop   /Selects between Position Feedback and Open Loop �                       ECS|Throttle1|Chan2ControlMode   Position Feedback|Open Loop   /Selects between Position Feedback and Open Loop �                      ECS|Throttle1|HP-EGRDC2Pos   V|%     �     	  @@ ����  X @@ ����  Y 
 P        ?   @��       B�            ECS|Throttle1|HP-EGRPosCal   V|%     �     	  @@ ����  X @@ ����  Y 
 P        ?   @��       B�            #ECS|Throttle1|Throttle1ModuleEnable   Enabled|Disabled   Enable Throttle �     !              ECS|Throttle1|Throttle1_Analog1   V     �     	    ??�            ECS|Throttle1|Throttle1_Analog2   V     �     	    ?p             'ECS|Throttle1|Throttle1_BattCompEnable1   |     �     !             'ECS|Throttle1|Throttle1_BattCompEnable2   |     �     !               ECS|Throttle1|Throttle1_BattNom1   V     �     	    A\��           ECS|Throttle1|Throttle1_BattNom2   V     �     	    A\��          ECS|Throttle1|Throttle1_Battery   V     �     	    A[�            &ECS|Throttle1|Throttle1_ControlEnable1   Enabled|Disabled   Enable Throttle �     !              &ECS|Throttle1|Throttle1_ControlEnable2   Enabled|Disabled   Enable Throttle �     !              ECS|Throttle1|Throttle1_Fault1    Fault|No Fault     �     !               ECS|Throttle1|Throttle1_Fault2    Fault|No Fault     �     !                ECS|Throttle1|Throttle1_I Sense1   A     �     	    =s�            ECS|Throttle1|Throttle1_I Sense2   A     �     	    =X�+           ECS|Throttle1|Throttle1_KRneg1   V/deg     �     	    ?333          ECS|Throttle1|Throttle1_KRneg2   V/deg     �     	    ?333          ECS|Throttle1|Throttle1_KRpos1   V/deg     �     	    ?             ECS|Throttle1|Throttle1_KRpos2   V/deg     �     	    ?333          (ECS|Throttle1|Throttle1_MotorResistance1   Ohms     �     	    @             (ECS|Throttle1|Throttle1_MotorResistance2   Ohms     �     	    @             ECS|Throttle1|Throttle1_Present   Present|Missing     �     !               ECS|Throttle1|Throttle1_TDneg1   s     �     	    <#�
          ECS|Throttle1|Throttle1_TDneg2   s     �     	    <#�
          ECS|Throttle1|Throttle1_TDpos1   s     �     	    <#�
          ECS|Throttle1|Throttle1_TDpos2   s     �     	    <#�
          ECS|Throttle1|Throttle1_TIneg1   s     �     	    >��          ECS|Throttle1|Throttle1_TIneg2   s     �     	    >��          ECS|Throttle1|Throttle1_TIpos1   s     �     	    >��          ECS|Throttle1|Throttle1_TIpos2   s     �     	    >��          ECS|Throttle1|Throttle1_TLag1   s     �     	    =L��          ECS|Throttle1|Throttle1_TLag2   s     �     	    =L��          ECS|Throttle1|Throttle1_TLead1   s     �     	                  ECS|Throttle1|Throttle1_TLead2   s     �     	                  #ECS|Throttle1|Throttle1_Temperature   C     �     	    A�Yl            ECS|Throttle1|Throttle1_ThetaLH1   deg     �     	                   ECS|Throttle1|Throttle1_ThetaLH2   deg     �     	                  +ECS|Throttle1|Throttle1_ThetaLHErrorThresh1   deg     �     	    >���          +ECS|Throttle1|Throttle1_ThetaLHErrorThresh2   deg     �     	    >���          ECS|Throttle1|Throttle1_ULH1   V     �     	    ?�            ECS|Throttle1|Throttle1_ULH2   V     �     	    ?�            ECS|Throttle1|Throttle1_ULHLag1   s     �     	    =u          ECS|Throttle1|Throttle1_ULHLag2   s     �     	    =u          ECS|Throttle1|Throttle1_US1   V     �     	    ?             ECS|Throttle1|Throttle1_US2   V     �     	    ?             ECS|Throttle1|Throttle1_USLag1   s     �     	    >��          ECS|Throttle1|Throttle1_USLag2   s     �     	    >��          ECS|Throttle|DesThrottleAngle   deg   -Desired Throttle Angle before manual settings �     	                   ECS|Throttle|DesThrottleDC   %   2Desired Throttle Duty Cycle before manual settings �     	    B��           #ECS|Throttle|DieselThrottleCalTable   mm3/cyc|rpm|%Open   Throttle Calibration Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B  B  B      D/  D;� DT� Dz  D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  ECS|Throttle|ManualThrottleAngle   deg   Manual Throttle Angle �     	    A�            &ECS|Throttle|ManualThrottleAngleEnable   Manual|Automatic   Enable Manual Throttle Angle �     !             ECS|Throttle|ManualThrottleDC   %   Manual Throttle Duty Cycle �     	    @�            #ECS|Throttle|ManualThrottleDCEnable   Manual|Automatic   !Enable Manual Throttle Duty Cycle �     !              !ECS|Throttle|Pedal2Throttle_Table   %|% Open     �     	  @@ ����  X @@ ����  Y 
 P            B�         B�            ECS|Throttle|Thr_Angle-DC_Table   %Open|%   Throttle Calibration Table �     	  @@ ����  X @@ ����  Y 
 P        @   B�33   @�  B�            ECS|Throttle|ThrottleAngle   %Open   Final Throttle Angle �     	    A�             ECS|Throttle|ThrottleDC   %   Final Throttle Duty Cycle �     	    B��           ECS|Throttle|ThrottlePosCal   V|%     �     	  @@ ����  X @@ ����  Y 
 P        ?   @��       B�            ECS|Torque|DesFuel   mm3/cyc   .Desired Fuel from table before manual override �     	                   ECS|Torque|DesFuelTable   Nm|RPM|mm3/cyc   Desired Fuel Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             @�  A�  BH  B�  B�  B�  C  C/  CH  Cz  C�  C�  C�  C�  C�     Cz  C�  D;� Dz  D�@ D�� D�� D�  E� E@ E+� E;� EZ� Ez  E�� E�@                                                                       ?�Q�?�Q�?�
=?�z�?�33?���?��\?(��?
=q>��>���>Ǯ>��R>�33>�p�>�p�@�  @�  @���@���@�ff@�33@y��@l��@Vff@@  @333@&ff@ff@��@   @   A��A��A��A  A33@���@�ff@�  @�33@�ff@�33@�  @�  @�  @ə�@ə�Ax  Ax  Al  A`  AT  AH  AA��A;33A8��A6ffA0  A)��A!��A!��A1��A1��A�ffA�ffA���A�33A���A�  A�33A�ffA���A���A|  AvffAk33Ak33Ay��Ay��A�ffA�ffA���A�33A���A�  A���A���A�ffA�33A���A�ffA���A���A�  A�  B  B  B  B  A�  A���A�33A�  A�33A�ffA�ffA�ffA�ffA�33A�ffA�ffBfffBfffBK��B0��B  B33A���A�  A�  A�  A�  A�  A�  A噚A�  A�  B�ffB�ffB�  B]33B6ffB  B  B33B  B��B��B
��B  B��B
  B
  B�  B�  B�ffB�33B�  BX��B@  B5��B3��B1��B133B0��B.  B2  B9��B9��B�33B�33B�  B�  B�� B�ffBp  B^ffB\  BY��BY  BXffB\ffBdffBnffBnffB�ffB�ffB�33B�33B�  B�33B�  B�ffB�  B�33B���B�  B�ffB���B���B���Bș�Bș�B�ffB�ffB�33B�33B���B���B�L�B���B��B�ffB�ffB�ffB�ffB�ffB���B���Bș�B�  B�ffB�  B�  B�  B��fBÙ�B��3B���B���B�  B�=qB���B�  B�  B���B���Bș�B�33B�33B�33B�  B�  B�  B�  B�  B�  B�  B�            ECS|Torque|DesTorque   Nm   "Desired Torque setpoint from table �     	                   ECS|Torque|DesTorqueTable   %|RPM|Nm   Torque Calibration Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P         	    ?� �@�  AH  A�  B3��B�B���B�         C�  Dz  D�� D�  E@ E;� EZ� Ez  E�� E�@ E�� E�    	                                                                                                               B�ffA�  Ah  @�ff                                    C
  B�33B  A���AH  @�ff@���                        C>33C�fB���BH��A�  A�33AH  A33@ٙ�                C�&fCv�C_�fCF��C&  B뙚B�  B5��A�33AH              C�  C�� C�  C�  C�  C�� Ci  CM  C)  B�ffA�          C�@ C�@ C�@ C�@ C���C�� C�  C�  C�  Ct  B           C�@ C�@ C�@ C�@ Cʙ�C�� C�  C�  C�  C�  Bp                ECS|Trig|9411_DigInput       +Logic level of the associated digital input �            ?           ECS|Trig|Digital_DC_Array   %   &Measured duty cycles of digital inputs �     	   @ ����       
                                               	    ECS|Trig|Digital_Freq_Array   Hz   $Measured frequency of digital inputs �     	   @ ����       
                                               	    ECS|Trig|Digital_PW_Array   Hz   'Measured pulse widths of digital inputs �     	   @ ����       
                                               	    ECS|UEGO1|Battery   V   Module Battery Voltage �     	    B�=           ECS|UEGO1|EGO1 Enable   Enabled|Disabled   Enable �     !              ECS|UEGO1|EGO1_Sensor   V   EGO Sensor Voltage �     	    >�ff           ECS|UEGO1|EGO1_Status   #COLD SENSOR|FOULED SENSOR|RICH|LEAN   EGO Sensor Status �                        ECS|UEGO1|EGO2 Enable   Enabled|Disabled   Enable �     !              ECS|UEGO1|EGO2_Sensor   V   EGO Sensor Voltage �     	    >�ff           ECS|UEGO1|EGO2_Status   #COLD SENSOR|FOULED SENSOR|RICH|LEAN   EGO Sensor Status �                        ECS|UEGO1|EGO3 Enable   Enabled|Disabled   Enable �     !              ECS|UEGO1|EGO3_Sensor   V   EGO Sensor Voltage �     	    >�ff           ECS|UEGO1|EGO3_Status   #COLD SENSOR|FOULED SENSOR|RICH|LEAN   EGO Sensor Status �                        ECS|UEGO1|EGO4 Enable   Enabled|Disabled   Enable �     !              ECS|UEGO1|EGO4_Sensor   V   EGO Sensor Voltage �     	    >�ff           ECS|UEGO1|EGO4_Status   #COLD SENSOR|FOULED SENSOR|RICH|LEAN   EGO Sensor Status �                        ECS|UEGO1|Fuse_Status   FUSE OK|FUSE BLOWN     �                        ECS|UEGO1|Module Enable   Enabled|Disabled   Override Backpressure �     !             ECS|UEGO1|Module_Present   Present|Missing   UEGO Module Present �     !              ECS|UEGO1|UEGO1 Back Pressure   bar   Back Pressure �     	    ?���           ECS|UEGO1|UEGO1 Enable   Enabled|Disabled   Enable �     !             $ECS|UEGO1|UEGO1 Manual Back Pressure   bar   Manual Back Pressure �     	    ?���          &ECS|UEGO1|UEGO1 Override Back Pressure   Manual|Automatic   Override Backpressure �     !              ECS|UEGO1|UEGO1_AF_Ratio       Air Fuel Ratio �     	    Ak33           !ECS|UEGO1|UEGO1_Heater_Duty_Cycle   %   UEGO heater duty cycle �     	                   ECS|UEGO1|UEGO1_Heater_Fault   6NO FAULT|SHORT TO BATTERY|OPEN CIRCUIT|SHORT TO GROUND     �                        ECS|UEGO1|UEGO1_Hot   Hot|Cold   
Sensor Hot �     !               ECS|UEGO1|UEGO1_Ip   mA   UEGO Current �     	                   ECS|UEGO1|UEGO1_Lambda       Lambda �     	    ?�             ECS|UEGO1|UEGO1_Phi       Phi �     	    ?�             ECS|UEGO1|UEGO1_Sensor_Fault   NO FAULT|SHORT TO GND OR BATT     �                        ECS|UEGO1|UEGO1_Temp   C   UEGO Temperature �     	    C�             ECS|UEGO1|UEGO2 Back Pressure   bar   Back Pressure �     	    ?���           ECS|UEGO1|UEGO2 Enable   Enabled|Disabled   Enable �     !             $ECS|UEGO1|UEGO2 Manual Back Pressure   bar   Manual Back Pressure �     	    ?���          &ECS|UEGO1|UEGO2 Override Back Pressure   Manual|Automatic   Override Backpressure �     !              ECS|UEGO1|UEGO2_AF_Ratio       Air Fuel Ratio �     	    Ak33           !ECS|UEGO1|UEGO2_Heater_Duty_Cycle   %   UEGO heater duty cycle �     	                   ECS|UEGO1|UEGO2_Heater_Fault   6NO FAULT|SHORT TO BATTERY|OPEN CIRCUIT|SHORT TO GROUND     �                        ECS|UEGO1|UEGO2_Hot   Hot|Cold   
Sensor Hot �     !               ECS|UEGO1|UEGO2_Ip   mA   UEGO Current �     	                   ECS|UEGO1|UEGO2_Lambda       Lambda �     	    ?�             ECS|UEGO1|UEGO2_Phi       Phi �     	    ?�             ECS|UEGO1|UEGO2_Sensor_Fault   NO FAULT|SHORT TO GND OR BATT     �                        ECS|UEGO1|UEGO2_Temp   C   UEGO Temperature �     	    C�             ECS|VVT|Cam1Angle_VVTSetpoint   mm3/cyc|rpm|deg   VVT Cam 1 Calibration Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B  B  B      D/  D;� DT� Dz  D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ�           B�  B�  B�  B�  B�  B�  B�  B�  BL  B  Ap              B�  B�  B�  B�  B�  B�  B�  B�  BL  B  Ap              B�  B�  B�  B�  B�  B�  B�  Bw33B8��A���Ap              B�  B�  B�  B�  Bp  Bp  Bp  B^  B(  A�  Ap              B�  B�  B�  Bh  BC  BC  BC  B2�B  A�
=@�              Bp  Bp  Bp  BD  B  B  B  B  A�  A4                  BH  BH  BH  B  B  B  B  A�
=A�  A"{                B%  B%  B%  B  A�  A�  A�  A�  A�  A                  B  B  B  A�  A�  A�  A�  A���A\��@���                B  B  B  A�  Ap  Ap  Ap  AX  A  @�                  A�  A�  A�  A�  @�  @�  @�  @ə�@�ff@ff                A�  A�  A�  A8                                          Ap  Ap  Ap  @�                                          @�  @�  @�  @`                                                                                                                                                                ECS|VVT|Cam1_Capture_End   DBTDC   0End of angle-based capture window for cam signal �     	    �p            ECS|VVT|Cam1_Capture_Start   DBTDC   2Start of angle-based capture window for cam signal �     	    Bp            ECS|VVT|Cam1_RisingEdge   DBTDC   !Captured angle of rising cam edge �     	                   ECS|VVT|Cam2Angle_VVTSetpoint   mm3/cyc|rpm|deg   VVT Cam 1 Calibration Table �     	  @@ ����  X @@ ����  Y @@ ��������  Z  P             @�  @�  A   AH  Ap  A�  A�  A�  A�  A�  A�  B  B  B  B      D/  D;� DT� Dz  D�@ D�� D�� D�  E� E@ E+� E;� EK  EZ�           B�  B�  B�  B�  B�  B�  B�  B�  BL  B  Ap              B�  B�  B�  B�  B�  B�  B�  B�  BL  B  Ap              B�  B�  B�  B�  B�  B�  B�  Bw33B8��A���Ap              B�  B�  B�  B�  Bp  Bp  Bp  B^  B(  A�  Ap              B�  B�  B�  Bh  BC  BC  BC  B2�B  A�
=@�              Bp  Bp  Bp  BD  B  B  B  B  A�  A4                  BH  BH  BH  B  B  B  B  A�
=A�  A"{                B%  B%  B%  B  A�  A�  A�  A�  A�  A                  B  B  B  A�  A�  A�  A�  A���A\��@���                B  B  B  A�  Ap  Ap  Ap  AX  A  @�                  A�  A�  A�  A�  @�  @�  @�  @ə�@�ff@ff                A�  A�  A�  A8                                          Ap  Ap  Ap  @�                                          @�  @�  @�  @`                                                                                                                                                                ECS|VVT|Cam2_Capture_End   DBTDC   0End of angle-based capture window for cam signal �     	    �p            ECS|VVT|Cam2_Capture_Start   DBTDC   2Start of angle-based capture window for cam signal �     	    Bp            ECS|VVT|Cam2_RisingEdge   DBTDC   !Captured angle of rising cam edge �     	                   ECS|VVT|CamRE_TDC-Ref   'TDC1|TDC2|TDC3|TDC4|TDC5|TDC6|TDC7|TDC8   @Selects Top Dead Center reference associated with driver channel �                       ECS|VVT|VVTCam1_ControlEnable   |   Enables PWM control of IMV �     !              ECS|VVT|VVTCam1_Current   A   QEstimated current to IMV based on battery voltage and nominal solenoid resistance �     	                   ECS|VVT|VVTCam1_DC   %   Final IMV duty cycle �     	                   ECS|VVT|VVTCam1_Freq   Hz   &Operating Frequency of IMV PWM command �     	    C/            ECS|VVT|VVTCam1_Kc   %/bar   IMV PID proportional gain �     	    :�o          ECS|VVT|VVTCam1_Kp_Action   %   /Proportional contribution of IMV PID controller �     	                   ECS|VVT|VVTCam1_ManualDC   %   ?Value to override IMV PID final output when ManualOverride=TRUE �     	                  ECS|VVT|VVTCam1_ManualOverride   |   0Causes ManualDC to override IMV PID final output �     !              ECS|VVT|VVTCam1_MaxDC   %   XMaximum allowed duty cycle for IMV. This value is effective if lower than IMV_MaxDCCalc. �     	                  ECS|VVT|VVTCam1_MaxDCCalc   %   �Maximum allowed duty cycle for IMV based on battery voltage and nominal solenoid resistance to limit current to 3A for channel pair �     	                   ECS|VVT|VVTCam1_MinDC   %   "Minimum allowed duty cycle for IMV �     	                  ECS|VVT|VVTCam1_NomResistance   Ohms   "Nominal resistance of IMV solenoid �     	    @             ECS|VVT|VVTCam1_NonPIDFF   %   FDuty cycle feed forward for the IMV while doing PID control of the HPV �     	    A�            ECS|VVT|VVTCam1_PID   %   pIMV PID controller output added to IMVPIDFF. Result is directed to selected PFI LS channel duty cycle parameter. �     	                   ECS|VVT|VVTCam1_PIDEnable   |   Enables PWM control of IMV �     !              ECS|VVT|VVTCam1_PIDFF   %   3Duty cycle feed forward added to the IMV PID output �     	    A�            ECS|VVT|VVTCam1_PIDMax   %   ;IMV PID output maximum limit (before feed forward is added) �     	    A�            ECS|VVT|VVTCam1_PIDMin   %   ;IMV PID output minimum limit (before feed forward is added) �     	    ��            ECS|VVT|VVTCam1_Td   min   YDerivative time constant for IMV PID controller (higher = stronger action. 0 = disabled.) �     	                  ECS|VVT|VVTCam1_Td_Action   A   -Derivative contribution of IMV PID controller �     	                   ECS|VVT|VVTCam1_Ti   min   VIntegral time constant for IMV PID controller (lower = stronger action. 0 = disabled.) �     	                  ECS|VVT|VVTCam1_Ti_Action   %   +Integral contribution of IMV PID controller �     	                   ECS|VVT|VVTCam2_ControlEnable   |   Enables PWM control of IMV �     !              ECS|VVT|VVTCam2_Current   A   QEstimated current to IMV based on battery voltage and nominal solenoid resistance �     	                   ECS|VVT|VVTCam2_DC   %   Final IMV duty cycle �     	                   ECS|VVT|VVTCam2_Freq   Hz   &Operating Frequency of IMV PWM command �     	    C/            ECS|VVT|VVTCam2_Kc   %/bar   IMV PID proportional gain �     	    :�o          ECS|VVT|VVTCam2_Kp_Action   %   /Proportional contribution of IMV PID controller �     	                   ECS|VVT|VVTCam2_ManualDC   %   ?Value to override IMV PID final output when ManualOverride=TRUE �     	                  ECS|VVT|VVTCam2_ManualOverride   |   0Causes ManualDC to override IMV PID final output �     !              ECS|VVT|VVTCam2_MaxDC   %   XMaximum allowed duty cycle for IMV. This value is effective if lower than IMV_MaxDCCalc. �     	                  ECS|VVT|VVTCam2_MaxDCCalc   %   �Maximum allowed duty cycle for IMV based on battery voltage and nominal solenoid resistance to limit current to 3A for channel pair �     	                   ECS|VVT|VVTCam2_MinDC   %   "Minimum allowed duty cycle for IMV �     	                  ECS|VVT|VVTCam2_NomResistance   Ohms   "Nominal resistance of IMV solenoid �     	    @             ECS|VVT|VVTCam2_NonPIDFF   %   FDuty cycle feed forward for the IMV while doing PID control of the HPV �     	    A�            ECS|VVT|VVTCam2_PID   %   pIMV PID controller output added to IMVPIDFF. Result is directed to selected PFI LS channel duty cycle parameter. �     	                   ECS|VVT|VVTCam2_PIDEnable   |   Enables PWM control of IMV �     !              ECS|VVT|VVTCam2_PIDFF   %   3Duty cycle feed forward added to the IMV PID output �     	    A�            ECS|VVT|VVTCam2_PIDMax   %   ;IMV PID output maximum limit (before feed forward is added) �     	    A�            ECS|VVT|VVTCam2_PIDMin   %   ;IMV PID output minimum limit (before feed forward is added) �     	    ��            ECS|VVT|VVTCam2_Td   min   YDerivative time constant for IMV PID controller (higher = stronger action. 0 = disabled.) �     	                  ECS|VVT|VVTCam2_Td_Action   A   -Derivative contribution of IMV PID controller �     	                   ECS|VVT|VVTCam2_Ti   min   VIntegral time constant for IMV PID controller (lower = stronger action. 0 = disabled.) �     	                  ECS|VVT|VVTCam2_Ti_Action   %   +Integral contribution of IMV PID controller �     	                   ECS|WG|WGEnable   |     �     !              ECS|WG|WGFreq         �     	               